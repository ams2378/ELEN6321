.subckt sbox a7 a6 a5 a4 a3 a2 a1 a0 d7 d6 d5 d4 d3 d2 d1 d0 gnd vdd
x1OR2X1TS n3202 n3556 n3563 gnd vdd OR2X1TS
x2NOR2X1TS n2617 n2716 n2819 gnd vdd NOR2X1TS
x3NAND2X1TS n2618 n2851 n2744 gnd vdd NAND2X1TS
x4NAND2X1TS n2619 n3391 n2618 gnd vdd NAND2X1TS
x5NOR2X1TS n2620 n2617 n2619 gnd vdd NOR2X1TS
x6NAND2X1TS n2621 n3018 n2620 gnd vdd NAND2X1TS
x7NOR2X1TS n2622 n2838 n2774 gnd vdd NOR2X1TS
x8NOR2X1TS n2623 n2771 n2768 gnd vdd NOR2X1TS
x9NOR2X1TS n2624 n3222 n2704 gnd vdd NOR2X1TS
x10NOR2X1TS n2625 n2782 n2815 gnd vdd NOR2X1TS
x11NOR2X1TS n2626 n2622 n2623 gnd vdd NOR2X1TS
x12NOR2X1TS n2627 n2624 n2625 gnd vdd NOR2X1TS
x13NAND2X1TS n2628 n2626 n2627 gnd vdd NAND2X1TS
x14NOR2X1TS n2629 n3357 n3358 gnd vdd NOR2X1TS
x15NAND2X1TS n2630 n3085 n3356 gnd vdd NAND2X1TS
x16NAND2X1TS n2631 n2629 n2630 gnd vdd NAND2X1TS
x17NOR2X1TS n2632 n2628 n2631 gnd vdd NOR2X1TS
x18NAND2X1TS n2633 n3017 n2632 gnd vdd NAND2X1TS
x19NOR2X1TS n2634 n2621 n2633 gnd vdd NOR2X1TS
x20NAND2X1TS n2635 n2965 n2634 gnd vdd NAND2X1TS
x21NOR2BX1TS n3060 n2955 n2635 gnd vdd NOR2BX1TS
x22NAND2X1TS n2636 n2877 n2784 gnd vdd NAND2X1TS
x23NAND2X1TS n2637 n3391 n2636 gnd vdd NAND2X1TS
x24NOR2X1TS n2638 n3462 n3463 gnd vdd NOR2X1TS
x25NOR2X1TS n2639 n2894 n3461 gnd vdd NOR2X1TS
x26NAND2X1TS n2640 n2871 n2639 gnd vdd NAND2X1TS
x27NAND2X1TS n2641 n2638 n2640 gnd vdd NAND2X1TS
x28NAND2X1TS n2642 n3004 n3458 gnd vdd NAND2X1TS
x29NAND2X1TS n2643 n3114 n2642 gnd vdd NAND2X1TS
x30NOR2X1TS n2644 n2831 n2982 gnd vdd NOR2X1TS
x31NOR2X1TS n2645 n2788 n2990 gnd vdd NOR2X1TS
x32NOR2X1TS n2646 n2641 n2643 gnd vdd NOR2X1TS
x33NOR2X1TS n2647 n2644 n2645 gnd vdd NOR2X1TS
x34NAND2X1TS n2648 n2646 n2647 gnd vdd NAND2X1TS
x35NOR2X1TS n2649 n2794 n3095 gnd vdd NOR2X1TS
x36NOR2X1TS n2650 n2637 n2648 gnd vdd NOR2X1TS
x37NOR2X1TS n2651 n3176 n2649 gnd vdd NOR2X1TS
x38NAND2X1TS n2652 n2650 n2651 gnd vdd NAND2X1TS
x39NAND2BX1TS n2653 n2652 n3248 gnd vdd NAND2BX1TS
x40NOR2X1TS n2654 n3053 n2653 gnd vdd NOR2X1TS
x41NAND2X1TS d0 n3164 n2654 gnd vdd NAND2X1TS
x42AND2X1TS n3141 n3428 n3500 gnd vdd AND2X1TS
x43NOR2BX1TS n2655 n3248 n3165 gnd vdd NOR2BX1TS
x44NAND2X1TS n2656 n2787 n2778 gnd vdd NAND2X1TS
x45NAND2X1TS n2657 n3115 n2737 gnd vdd NAND2X1TS
x46NAND2X1TS n2658 n2656 n2657 gnd vdd NAND2X1TS
x47NAND2X1TS n2659 n3220 n3219 gnd vdd NAND2X1TS
x48NOR2X1TS n2660 n3223 n3224 gnd vdd NOR2X1TS
x49NAND2X1TS n2661 n2745 n3221 gnd vdd NAND2X1TS
x50NAND2X1TS n2662 n2660 n2661 gnd vdd NAND2X1TS
x51NOR2X1TS n2663 n2833 n2807 gnd vdd NOR2X1TS
x52AND2X1TS n2664 n2846 n2748 gnd vdd AND2X1TS
x53NOR2X1TS n2665 n2659 n2662 gnd vdd NOR2X1TS
x54NOR2X1TS n2666 n2663 n2664 gnd vdd NOR2X1TS
x55NAND2X1TS n2667 n2665 n2666 gnd vdd NAND2X1TS
x56NOR2X1TS n2668 n2658 n2667 gnd vdd NOR2X1TS
x57NAND2X1TS n2669 n3031 n2668 gnd vdd NAND2X1TS
x58NOR2X1TS n2670 n2669 n3179 gnd vdd NOR2X1TS
x59NOR2X1TS n2671 n3196 n3203 gnd vdd NOR2X1TS
x60NAND2X1TS n2672 n2670 n2671 gnd vdd NAND2X1TS
x61NOR2X1TS n2673 n3247 n2672 gnd vdd NOR2X1TS
x62NAND2X1TS d2 n2655 n2673 gnd vdd NAND2X1TS
x63NOR2X1TS n2674 n2840 n3171 gnd vdd NOR2X1TS
x64NOR2X1TS n2675 n2830 n2712 gnd vdd NOR2X1TS
x65NOR2X1TS n2676 n2674 n2675 gnd vdd NOR2X1TS
x66NAND2X1TS n2677 n2851 n2779 gnd vdd NAND2X1TS
x67NAND2X1TS n2678 n2676 n2677 gnd vdd NAND2X1TS
x68NAND2X1TS n2679 n2726 n3170 gnd vdd NAND2X1TS
x69NAND2X1TS n2680 n2785 n3166 gnd vdd NAND2X1TS
x70NAND2X1TS n2681 n2679 n2680 gnd vdd NAND2X1TS
x71NOR2BX1TS n2682 n2849 n3167 gnd vdd NOR2BX1TS
x72NOR2X1TS n2683 n2682 n2681 gnd vdd NOR2X1TS
x73NAND2X1TS n2684 n2933 n3168 gnd vdd NAND2X1TS
x74NAND2X1TS n2685 n2683 n2684 gnd vdd NAND2X1TS
x75NOR2X1TS n2686 n2719 n2761 gnd vdd NOR2X1TS
x76NOR2X1TS n2687 n3172 n2686 gnd vdd NOR2X1TS
x77NAND2X1TS n2688 n3070 n2687 gnd vdd NAND2X1TS
x78NOR2X1TS n2689 n2678 n2685 gnd vdd NOR2X1TS
x79NOR2X1TS n2690 n2688 n3165 gnd vdd NOR2X1TS
x80NAND2X1TS n2691 n2689 n2690 gnd vdd NAND2X1TS
x81NOR2X1TS n2692 n3028 n2691 gnd vdd NOR2X1TS
x82NAND2X1TS d3 n3164 n2692 gnd vdd NAND2X1TS
x83AND2X2TS n2693 n3500 n3555 gnd vdd AND2X2TS
x84AND2X2TS n2694 n2706 n3555 gnd vdd AND2X2TS
x85AND2X2TS n2695 n3500 n3460 gnd vdd AND2X2TS
x86AND2X2TS n2696 n2913 n3446 gnd vdd AND2X2TS
x87OR2X2TS n2697 n3568 n3569 gnd vdd OR2X2TS
x88AND2X2TS n2698 n3446 n3562 gnd vdd AND2X2TS
x89AND2X2TS n2699 n2903 n3304 gnd vdd AND2X2TS
x90AND2X2TS n2700 n3499 n3459 gnd vdd AND2X2TS
x91AND2X2TS n2701 n3370 n3466 gnd vdd AND2X2TS
x92OR2X2TS n2702 n2863 n2857 gnd vdd OR2X2TS
x93NAND2X1TS n2703 n2905 n2893 gnd vdd NAND2X1TS
x94INVXLTS n2704 n2994 gnd vdd INVXLTS
x95INVXLTS n2705 n2994 gnd vdd INVXLTS
x96INVXLTS n2706 n2703 gnd vdd INVXLTS
x97INVXLTS n2707 n2703 gnd vdd INVXLTS
x98INVXLTS n2708 n3460 gnd vdd INVXLTS
x99INVXLTS n2709 n2708 gnd vdd INVXLTS
x100INVXLTS n2710 n2933 gnd vdd INVXLTS
x101INVXLTS n2711 n2702 gnd vdd INVXLTS
x102INVXLTS n2712 n2702 gnd vdd INVXLTS
x103INVXLTS n2713 n3096 gnd vdd INVXLTS
x104INVXLTS n2714 n3096 gnd vdd INVXLTS
x105INVXLTS n2715 n2939 gnd vdd INVXLTS
x106INVXLTS n2716 n2939 gnd vdd INVXLTS
x107INVXLTS n2717 n3131 gnd vdd INVXLTS
x108INVXLTS n2718 n3131 gnd vdd INVXLTS
x109INVXLTS n2719 n2925 gnd vdd INVXLTS
x110INVXLTS n2720 n2925 gnd vdd INVXLTS
x111INVXLTS n2721 n2975 gnd vdd INVXLTS
x112INVXLTS n2722 n2975 gnd vdd INVXLTS
x113INVXLTS n2723 n2700 gnd vdd INVXLTS
x114INVXLTS n2724 n2700 gnd vdd INVXLTS
x115INVXLTS n2725 n3202 gnd vdd INVXLTS
x116INVXLTS n2726 n3202 gnd vdd INVXLTS
x117INVXLTS n2727 n2935 gnd vdd INVXLTS
x118INVXLTS n2728 n2935 gnd vdd INVXLTS
x119INVXLTS n2729 n2697 gnd vdd INVXLTS
x120INVXLTS n2730 n2697 gnd vdd INVXLTS
x121INVXLTS n2731 n2699 gnd vdd INVXLTS
x122INVXLTS n2732 n2699 gnd vdd INVXLTS
x123INVXLTS n2733 n2698 gnd vdd INVXLTS
x124INVXLTS n2734 n2698 gnd vdd INVXLTS
x125INVXLTS n2735 n3161 gnd vdd INVXLTS
x126INVXLTS n2736 n3161 gnd vdd INVXLTS
x127INVXLTS n2737 n3080 gnd vdd INVXLTS
x128INVXLTS n2738 n3080 gnd vdd INVXLTS
x129INVXLTS n2739 n2701 gnd vdd INVXLTS
x130INVXLTS n2740 n2701 gnd vdd INVXLTS
x131INVXLTS n2741 n2945 gnd vdd INVXLTS
x132INVXLTS n2742 n2741 gnd vdd INVXLTS
x133INVXLTS n2743 n2741 gnd vdd INVXLTS
x134INVXLTS n2744 n2945 gnd vdd INVXLTS
x135INVXLTS n2745 n2945 gnd vdd INVXLTS
x136INVXLTS n2746 n3006 gnd vdd INVXLTS
x137INVXLTS n2747 n2746 gnd vdd INVXLTS
x138INVXLTS n2748 n2746 gnd vdd INVXLTS
x139INVXLTS n2749 n3023 gnd vdd INVXLTS
x140INVXLTS n2750 n2749 gnd vdd INVXLTS
x141INVXLTS n2751 n2988 gnd vdd INVXLTS
x142INVXLTS n2752 n2751 gnd vdd INVXLTS
x143INVXLTS n2753 n2751 gnd vdd INVXLTS
x144INVXLTS n2754 n3089 gnd vdd INVXLTS
x145INVXLTS n2756 n3089 gnd vdd INVXLTS
x146INVXLTS n2755 n3089 gnd vdd INVXLTS
x147INVXLTS n2757 n2928 gnd vdd INVXLTS
x148INVXLTS n2759 n2928 gnd vdd INVXLTS
x149INVXLTS n2758 n2928 gnd vdd INVXLTS
x150INVXLTS n2760 n2693 gnd vdd INVXLTS
x151INVXLTS n2762 n2693 gnd vdd INVXLTS
x152INVXLTS n2761 n2693 gnd vdd INVXLTS
x153INVXLTS n2763 n3125 gnd vdd INVXLTS
x154INVXLTS n2765 n3125 gnd vdd INVXLTS
x155INVXLTS n2764 n3125 gnd vdd INVXLTS
x156INVXLTS n2766 n2986 gnd vdd INVXLTS
x157INVXLTS n2768 n2986 gnd vdd INVXLTS
x158INVXLTS n2767 n2986 gnd vdd INVXLTS
x159INVXLTS n2769 n2760 gnd vdd INVXLTS
x160INVXLTS n2770 n2762 gnd vdd INVXLTS
x161INVXLTS n2772 n3051 gnd vdd INVXLTS
x162INVXLTS n2771 n3051 gnd vdd INVXLTS
x163INVXLTS n2773 n3013 gnd vdd INVXLTS
x164INVXLTS n2774 n2773 gnd vdd INVXLTS
x165INVXLTS n2776 n2773 gnd vdd INVXLTS
x166INVXLTS n2775 n2773 gnd vdd INVXLTS
x167INVXLTS n2777 n3085 gnd vdd INVXLTS
x168INVXLTS n2778 n2777 gnd vdd INVXLTS
x169INVXLTS n2779 n2777 gnd vdd INVXLTS
x170INVXLTS n2780 n3077 gnd vdd INVXLTS
x171INVXLTS n2782 n3077 gnd vdd INVXLTS
x172INVXLTS n2781 n3077 gnd vdd INVXLTS
x173INVXLTS n2783 n2791 gnd vdd INVXLTS
x174INVXLTS n2784 n2793 gnd vdd INVXLTS
x175INVXLTS n2785 n3013 gnd vdd INVXLTS
x176INVXLTS n2787 n3013 gnd vdd INVXLTS
x177INVXLTS n2786 n3013 gnd vdd INVXLTS
x178INVXLTS n2788 n2763 gnd vdd INVXLTS
x179INVXLTS n2790 n2765 gnd vdd INVXLTS
x180INVXLTS n2789 n2764 gnd vdd INVXLTS
x181INVXLTS n2791 n2695 gnd vdd INVXLTS
x182INVXLTS n2793 n2695 gnd vdd INVXLTS
x183INVXLTS n2792 n2695 gnd vdd INVXLTS
x184INVXLTS n2794 n2694 gnd vdd INVXLTS
x185INVXLTS n2796 n2694 gnd vdd INVXLTS
x186INVXLTS n2795 n2694 gnd vdd INVXLTS
x187INVXLTS n2798 n2988 gnd vdd INVXLTS
x188INVXLTS n2797 n2988 gnd vdd INVXLTS
x189INVXLTS n2799 n3015 gnd vdd INVXLTS
x190INVXLTS n2800 n2799 gnd vdd INVXLTS
x191INVXLTS n2801 n2799 gnd vdd INVXLTS
x192INVXLTS n2802 n3141 gnd vdd INVXLTS
x193INVXLTS n2804 n3141 gnd vdd INVXLTS
x194INVXLTS n2803 n3141 gnd vdd INVXLTS
x195INVXLTS n2805 n2946 gnd vdd INVXLTS
x196INVXLTS n2807 n2946 gnd vdd INVXLTS
x197INVXLTS n2806 n2946 gnd vdd INVXLTS
x198INVXLTS n2808 n2699 gnd vdd INVXLTS
x199INVXLTS n2809 n2808 gnd vdd INVXLTS
x200INVXLTS n2811 n2808 gnd vdd INVXLTS
x201INVXLTS n2810 n2808 gnd vdd INVXLTS
x202INVXLTS n2812 n3096 gnd vdd INVXLTS
x203INVXLTS n2813 n2812 gnd vdd INVXLTS
x204INVXLTS n2815 n2812 gnd vdd INVXLTS
x205INVXLTS n2814 n2812 gnd vdd INVXLTS
x206INVXLTS n2816 n2796 gnd vdd INVXLTS
x207INVXLTS n2817 n2794 gnd vdd INVXLTS
x208INVXLTS n2818 n3131 gnd vdd INVXLTS
x209INVXLTS n2819 n2818 gnd vdd INVXLTS
x210INVXLTS n2821 n2818 gnd vdd INVXLTS
x211INVXLTS n2820 n2818 gnd vdd INVXLTS
x212INVXLTS n2822 n2696 gnd vdd INVXLTS
x213INVXLTS n2824 n2696 gnd vdd INVXLTS
x214INVXLTS n2823 n2696 gnd vdd INVXLTS
x215INVXLTS n2825 n3080 gnd vdd INVXLTS
x216INVXLTS n2826 n2825 gnd vdd INVXLTS
x217INVXLTS n2828 n2825 gnd vdd INVXLTS
x218INVXLTS n2827 n2825 gnd vdd INVXLTS
x219INVXLTS n2829 n2755 gnd vdd INVXLTS
x220INVXLTS n2830 n2756 gnd vdd INVXLTS
x221INVXLTS n2831 n2754 gnd vdd INVXLTS
x222INVXLTS n2832 n3202 gnd vdd INVXLTS
x223INVXLTS n2835 n2832 gnd vdd INVXLTS
x224INVXLTS n2833 n2832 gnd vdd INVXLTS
x225INVXLTS n2834 n2832 gnd vdd INVXLTS
x226INVXLTS n2836 n2954 gnd vdd INVXLTS
x227INVXLTS n2837 n2836 gnd vdd INVXLTS
x228INVXLTS n2838 n2836 gnd vdd INVXLTS
x229INVXLTS n2839 n2836 gnd vdd INVXLTS
x230INVXLTS n2840 n3051 gnd vdd INVXLTS
x231INVXLTS n2841 n2840 gnd vdd INVXLTS
x232INVXLTS n2842 n2840 gnd vdd INVXLTS
x233INVXLTS n2843 n2700 gnd vdd INVXLTS
x234INVXLTS n2844 n2843 gnd vdd INVXLTS
x235INVXLTS n2846 n2843 gnd vdd INVXLTS
x236INVXLTS n2845 n2843 gnd vdd INVXLTS
x237INVXLTS n2847 n2946 gnd vdd INVXLTS
x238INVXLTS n2848 n2847 gnd vdd INVXLTS
x239INVXLTS n2849 n2847 gnd vdd INVXLTS
x240INVXLTS n2850 n3141 gnd vdd INVXLTS
x241INVXLTS n2851 n2850 gnd vdd INVXLTS
x242INVXLTS n2852 n2850 gnd vdd INVXLTS
x243INVXLTS n2853 n3161 gnd vdd INVXLTS
x244INVXLTS n2854 n2853 gnd vdd INVXLTS
x245INVXLTS n2855 n2853 gnd vdd INVXLTS
x246INVXLTS n2856 n2939 gnd vdd INVXLTS
x247INVXLTS n2857 n2856 gnd vdd INVXLTS
x248INVXLTS n2858 n2856 gnd vdd INVXLTS
x249INVXLTS n2859 n2767 gnd vdd INVXLTS
x250INVXLTS n2860 n2766 gnd vdd INVXLTS
x251INVXLTS n2861 n2933 gnd vdd INVXLTS
x252INVXLTS n2862 n2861 gnd vdd INVXLTS
x253INVXLTS n2863 n2861 gnd vdd INVXLTS
x254INVXLTS n2864 n3077 gnd vdd INVXLTS
x255INVXLTS n2865 n2864 gnd vdd INVXLTS
x256INVXLTS n2867 n2864 gnd vdd INVXLTS
x257INVXLTS n2866 n2864 gnd vdd INVXLTS
x258INVXLTS n2868 n2975 gnd vdd INVXLTS
x259INVXLTS n2869 n2868 gnd vdd INVXLTS
x260INVXLTS n2871 n2868 gnd vdd INVXLTS
x261INVXLTS n2870 n2868 gnd vdd INVXLTS
x262INVXLTS n2872 n2994 gnd vdd INVXLTS
x263INVXLTS n2873 n2872 gnd vdd INVXLTS
x264INVXLTS n2874 n2872 gnd vdd INVXLTS
x265INVXLTS n2875 n2872 gnd vdd INVXLTS
x266INVXLTS n2876 n2928 gnd vdd INVXLTS
x267INVXLTS n2877 n2876 gnd vdd INVXLTS
x268INVXLTS n2878 n2876 gnd vdd INVXLTS
x269INVXLTS n2879 n2876 gnd vdd INVXLTS
x270INVXLTS n2880 n2925 gnd vdd INVXLTS
x271INVXLTS n2881 n2880 gnd vdd INVXLTS
x272INVXLTS n2882 n2880 gnd vdd INVXLTS
x273INVXLTS n2883 n2880 gnd vdd INVXLTS
x274INVXLTS n2884 n2935 gnd vdd INVXLTS
x275INVXLTS n2885 n2884 gnd vdd INVXLTS
x276INVXLTS n2888 n2884 gnd vdd INVXLTS
x277INVXLTS n2886 n2884 gnd vdd INVXLTS
x278INVXLTS n2887 n2884 gnd vdd INVXLTS
x279INVXLTS n2889 a2 gnd vdd INVXLTS
x280INVXLTS n2890 n2889 gnd vdd INVXLTS
x281INVXLTS n2891 n2889 gnd vdd INVXLTS
x282INVXLTS n2892 a7 gnd vdd INVXLTS
x283INVXLTS n2893 n2892 gnd vdd INVXLTS
x284INVXLTS n2894 n2892 gnd vdd INVXLTS
x285INVXLTS n2895 a6 gnd vdd INVXLTS
x286INVXLTS n2896 n2895 gnd vdd INVXLTS
x287INVXLTS n2897 n2895 gnd vdd INVXLTS
x288INVXLTS n2898 a3 gnd vdd INVXLTS
x289INVXLTS n2899 n2898 gnd vdd INVXLTS
x290INVXLTS n2900 n2898 gnd vdd INVXLTS
x291INVXLTS n2901 a0 gnd vdd INVXLTS
x292INVXLTS n2902 n2901 gnd vdd INVXLTS
x293INVXLTS n2903 n2901 gnd vdd INVXLTS
x294INVXLTS n2904 a5 gnd vdd INVXLTS
x295INVXLTS n2905 n2904 gnd vdd INVXLTS
x296INVXLTS n2906 n2904 gnd vdd INVXLTS
x297INVXLTS n2907 a4 gnd vdd INVXLTS
x298INVXLTS n2908 n2907 gnd vdd INVXLTS
x299INVXLTS n2909 n2907 gnd vdd INVXLTS
x300INVXLTS n2910 a1 gnd vdd INVXLTS
x301INVXLTS n2911 n2910 gnd vdd INVXLTS
x302INVXLTS n2913 n2910 gnd vdd INVXLTS
x303INVXLTS n2912 n2910 gnd vdd INVXLTS
x304AND2XLTS n2718 n3464 n3463 gnd vdd AND2XLTS
x305NOR2XLTS n3462 n2736 n3465 gnd vdd NOR2XLTS
x306NOR2XLTS n2962 n2963 n2964 gnd vdd NOR2XLTS
x307NOR2XLTS n2966 n2967 n2968 gnd vdd NOR2XLTS
x308NOR2XLTS n2970 n2971 n2972 gnd vdd NOR2XLTS
x309NOR2XLTS n2971 n2977 n2734 gnd vdd NOR2XLTS
x310NOR2XLTS n2969 n2978 n2979 gnd vdd NOR2XLTS
x311NOR2XLTS n2990 n2750 n2745 gnd vdd NOR2XLTS
x312NOR2XLTS n2961 n2917 n2991 gnd vdd NOR2XLTS
x313NOR2XLTS n3027 n3028 n3029 gnd vdd NOR2XLTS
x314NOR2XLTS n3030 n3032 n3033 gnd vdd NOR2XLTS
x315NOR2XLTS n3035 n3036 n3037 gnd vdd NOR2XLTS
x316NOR2XLTS n3037 n2734 n2772 gnd vdd NOR2XLTS
x317NOR2XLTS n3034 n3038 n3039 gnd vdd NOR2XLTS
x318NOR2XLTS n3039 n2711 n2735 gnd vdd NOR2XLTS
x319NOR2XLTS n3038 n3040 n2805 gnd vdd NOR2XLTS
x320NOR2XLTS n3042 n3043 n3044 gnd vdd NOR2XLTS
x321AND2XLTS n2846 n2976 n3044 gnd vdd AND2XLTS
x322NOR2XLTS n3046 n2891 n2913 gnd vdd NOR2XLTS
x323NOR2XLTS n3043 n3047 n2710 gnd vdd NOR2XLTS
x324NOR2XLTS n3041 n3048 n3049 gnd vdd NOR2XLTS
x325NOR2XLTS n3049 n3050 n2739 gnd vdd NOR2XLTS
x326NOR2XLTS n3050 n2694 n2841 gnd vdd NOR2XLTS
x327NOR2XLTS n3048 n2839 n2947 gnd vdd NOR2XLTS
x328NOR2XLTS n3026 n3052 n3053 gnd vdd NOR2XLTS
x329OR2XLTS n3203 n3467 n3053 gnd vdd OR2XLTS
x330NOR2XLTS n3469 n3470 n3471 gnd vdd NOR2XLTS
x331NOR2XLTS n3470 n2831 n2824 gnd vdd NOR2XLTS
x332NOR2XLTS n3468 n3474 n3475 gnd vdd NOR2XLTS
x333NOR2XLTS n3479 n3483 n3484 gnd vdd NOR2XLTS
x334NOR2XLTS n3484 n3485 n2821 gnd vdd NOR2XLTS
x335NOR2XLTS n3485 n2858 n2878 gnd vdd NOR2XLTS
x336NOR2XLTS n3483 n3486 n2760 gnd vdd NOR2XLTS
x337NOR2XLTS n3486 n2867 n3446 gnd vdd NOR2XLTS
x338NOR2XLTS n3055 n3056 n3057 gnd vdd NOR2XLTS
x339NOR2XLTS n3056 n2804 n2758 gnd vdd NOR2XLTS
x340NOR2XLTS n3054 n3058 n3059 gnd vdd NOR2XLTS
x341NOR2XLTS n3061 n2963 n3062 gnd vdd NOR2XLTS
x342NOR2XLTS n3066 n3067 n3068 gnd vdd NOR2XLTS
x343NOR2XLTS n3067 n2837 n2806 gnd vdd NOR2XLTS
x344NOR2XLTS n3063 n3098 n3099 gnd vdd NOR2XLTS
x345NOR2XLTS n3106 n3107 n3108 gnd vdd NOR2XLTS
x346NOR2XLTS n3108 n3109 n2781 gnd vdd NOR2XLTS
x347NOR2XLTS n3107 n3110 n2804 gnd vdd NOR2XLTS
x348NOR2XLTS n3105 n3111 n3112 gnd vdd NOR2XLTS
x349NOR2XLTS n3111 n2719 n2732 gnd vdd NOR2XLTS
x350OR2XLTS n2953 n3116 n2963 gnd vdd OR2XLTS
x351NOR2XLTS n3118 n3119 n3120 gnd vdd NOR2XLTS
x352NOR2XLTS n3122 n3123 n3124 gnd vdd NOR2XLTS
x353NOR2XLTS n3124 n2705 n2790 gnd vdd NOR2XLTS
x354NOR2XLTS n3121 n3126 n3127 gnd vdd NOR2XLTS
x355NOR2XLTS n3126 n3133 n2735 gnd vdd NOR2XLTS
x356NOR2XLTS n3133 n2888 n3134 gnd vdd NOR2XLTS
x357NOR2XLTS n3119 n3135 n2815 gnd vdd NOR2XLTS
x358NOR2XLTS n3135 n3023 n3136 gnd vdd NOR2XLTS
x359NOR2XLTS n3117 n3137 n3138 gnd vdd NOR2XLTS
x360NOR2XLTS n2915 n2916 n2917 gnd vdd NOR2XLTS
x361NOR2XLTS n2996 n2997 n2998 gnd vdd NOR2XLTS
x362NOR2XLTS n3000 n3001 n3002 gnd vdd NOR2XLTS
x363NOR2XLTS n3002 n2977 n3003 gnd vdd NOR2XLTS
x364NOR2XLTS n3001 n3005 n2736 gnd vdd NOR2XLTS
x365NOR2XLTS n3005 n2881 n2748 gnd vdd NOR2XLTS
x366NOR2XLTS n2999 n3007 n3008 gnd vdd NOR2XLTS
x367NOR2XLTS n3009 n3011 n3012 gnd vdd NOR2XLTS
x368NOR2XLTS n3012 n2776 n2743 gnd vdd NOR2XLTS
x369NOR2XLTS n3011 n3014 n2801 gnd vdd NOR2XLTS
x370NOR2XLTS n3007 n3016 n2822 gnd vdd NOR2XLTS
x371NOR2XLTS n2995 n3019 n3020 gnd vdd NOR2XLTS
x372NOR2XLTS n3021 n3024 n3025 gnd vdd NOR2XLTS
x373NOR2XLTS n3025 n2759 n2771 gnd vdd NOR2XLTS
x374NOR2XLTS n3024 n2954 n2724 gnd vdd NOR2XLTS
x375NOR2XLTS n2919 n2920 n2921 gnd vdd NOR2XLTS
x376NOR2XLTS n2918 n2929 n2930 gnd vdd NOR2XLTS
x377NOR2XLTS n2937 n2942 n2943 gnd vdd NOR2XLTS
x378NOR2XLTS n2943 n2944 n2743 gnd vdd NOR2XLTS
x379NOR2XLTS n2944 n2763 n2848 gnd vdd NOR2XLTS
x380NOR2XLTS n2942 n2722 n2947 gnd vdd NOR2XLTS
x381NOR2XLTS n2914 n2948 n2949 gnd vdd NOR2XLTS
x382NOR2XLTS n2951 n3081 n3082 gnd vdd NOR2XLTS
x383NOR2XLTS n3083 n3086 n3087 gnd vdd NOR2XLTS
x384NOR2XLTS n3086 n3088 n2829 gnd vdd NOR2XLTS
x385NOR2XLTS n3090 n3093 n3094 gnd vdd NOR2XLTS
x386NOR2XLTS n3094 n3095 n2813 gnd vdd NOR2XLTS
x387NOR2XLTS n3095 n2778 n2869 gnd vdd NOR2XLTS
x388NOR2XLTS n3093 n3016 n2740 gnd vdd NOR2XLTS
x389NOR2XLTS n3016 n2816 n2784 gnd vdd NOR2XLTS
x390NOR2XLTS n2950 n2952 n2953 gnd vdd NOR2XLTS
x391NOR2XLTS n3145 n3146 n3147 gnd vdd NOR2XLTS
x392NOR2XLTS n3146 n3151 n2803 gnd vdd NOR2XLTS
x393NOR2XLTS n3144 n3152 n3153 gnd vdd NOR2XLTS
x394NOR2XLTS n3158 n2873 n2859 gnd vdd NOR2XLTS
x395NOR2XLTS n2982 n2750 n2863 gnd vdd NOR2XLTS
x396NOR2XLTS n2952 n2838 n2802 gnd vdd NOR2XLTS
x397NOR2XLTS n2956 n2957 n2958 gnd vdd NOR2XLTS
x398NOR2XLTS n2959 n3071 n3072 gnd vdd NOR2XLTS
x399NOR2XLTS n3075 n3078 n3079 gnd vdd NOR2XLTS
x400NOR2XLTS n3079 n2715 n2776 gnd vdd NOR2XLTS
x401NOR2XLTS n3078 n2757 n2826 gnd vdd NOR2XLTS
x402NOR2XLTS n3164 n3247 n3508 gnd vdd NOR2XLTS
x403OR2XLTS n3057 n3509 n3508 gnd vdd OR2XLTS
x404NOR2XLTS n3511 n3512 n3513 gnd vdd NOR2XLTS
x405NOR2XLTS n3514 n3516 n3517 gnd vdd NOR2XLTS
x406NOR2XLTS n3517 n3187 n2772 gnd vdd NOR2XLTS
x407NOR2XLTS n3516 n3518 n2768 gnd vdd NOR2XLTS
x408NOR2XLTS n3518 n2842 n2786 gnd vdd NOR2XLTS
x409NOR2XLTS n3512 n3218 n2752 gnd vdd NOR2XLTS
x410NOR2XLTS n3510 n3519 n3520 gnd vdd NOR2XLTS
x411INVXLTS n3458 n3222 gnd vdd INVXLTS
x412NOR2XLTS n3519 n3525 n2828 gnd vdd NOR2XLTS
x413NOR2XLTS n3525 n2702 n3136 gnd vdd NOR2XLTS
x414NOR2XLTS n3529 n3530 n3531 gnd vdd NOR2XLTS
x415NOR2XLTS n3531 n3151 n2736 gnd vdd NOR2XLTS
x416NOR2XLTS n3530 n3532 n2732 gnd vdd NOR2XLTS
x417NOR2XLTS n3532 n2875 n3424 gnd vdd NOR2XLTS
x418NOR2XLTS n3528 n3533 n3534 gnd vdd NOR2XLTS
x419NOR2XLTS n3535 n3536 n3537 gnd vdd NOR2XLTS
x420NOR2XLTS n3537 n2704 n2802 gnd vdd NOR2XLTS
x421NOR2XLTS n3536 n3169 n2834 gnd vdd NOR2XLTS
x422NOR2XLTS n3533 n3110 n2807 gnd vdd NOR2XLTS
x423INVXLTS n3110 n3136 gnd vdd INVXLTS
x424NOR2XLTS n3172 n2740 n2723 gnd vdd NOR2XLTS
x425NOR2XLTS n3174 n3175 n3176 gnd vdd NOR2XLTS
x426NOR2XLTS n3430 n3432 n3433 gnd vdd NOR2XLTS
x427NOR2XLTS n3178 n3179 n3180 gnd vdd NOR2XLTS
x428INVXLTS n3183 n3184 gnd vdd INVXLTS
x429NOR2XLTS n3181 n3185 n3186 gnd vdd NOR2XLTS
x430NOR2XLTS n3186 n3187 n2826 gnd vdd NOR2XLTS
x431NOR2XLTS n3187 n2873 n2877 gnd vdd NOR2XLTS
x432NOR2XLTS n3185 n3188 n2813 gnd vdd NOR2XLTS
x433NOR2XLTS n3188 n2887 n2879 gnd vdd NOR2XLTS
x434NOR2XLTS n3177 n3189 n3190 gnd vdd NOR2XLTS
x435NOR2XLTS n3189 n3195 n2705 gnd vdd NOR2XLTS
x436NOR2XLTS n3195 n2845 n2934 gnd vdd NOR2XLTS
x437NOR2XLTS n3173 n3196 n3197 gnd vdd NOR2XLTS
x438NOR2XLTS n3198 n3200 n3201 gnd vdd NOR2XLTS
x439NOR2XLTS n3201 n2819 n2835 gnd vdd NOR2XLTS
x440NOR2XLTS n3200 n2801 n2752 gnd vdd NOR2XLTS
x441NOR2XLTS n3205 n3087 n3206 gnd vdd NOR2XLTS
x442NOR2XLTS n3206 n2830 n2742 gnd vdd NOR2XLTS
x443NOR2XLTS n3087 n2760 n2721 gnd vdd NOR2XLTS
x444NOR2XLTS n3204 n3207 n3208 gnd vdd NOR2XLTS
x445NOR2XLTS n3208 n3015 n2827 gnd vdd NOR2XLTS
x446NOR2XLTS n3207 n3104 n2789 gnd vdd NOR2XLTS
x447NOR2XLTS n3210 n3211 n3212 gnd vdd NOR2XLTS
x448NOR2XLTS n3212 n3184 n2835 gnd vdd NOR2XLTS
x449NOR2XLTS n3184 n2764 n2841 gnd vdd NOR2XLTS
x450NOR2XLTS n3211 n3213 n2795 gnd vdd NOR2XLTS
x451NOR2XLTS n3213 n2933 n3166 gnd vdd NOR2XLTS
x452NOR2XLTS n3209 n3214 n3215 gnd vdd NOR2XLTS
x453NOR2XLTS n3214 n3218 n2807 gnd vdd NOR2XLTS
x454NOR2XLTS n3218 n2779 n2882 gnd vdd NOR2XLTS
x455NOR2XLTS n3488 n3364 n3489 gnd vdd NOR2XLTS
x456NOR2XLTS n3490 n3492 n3493 gnd vdd NOR2XLTS
x457NOR2XLTS n3493 n2829 n2722 gnd vdd NOR2XLTS
x458NOR2XLTS n3492 n2780 n2792 gnd vdd NOR2XLTS
x459NOR2XLTS n3487 n3494 n3495 gnd vdd NOR2XLTS
x460NOR2XLTS n3498 n2717 n2756 gnd vdd NOR2XLTS
x461NOR2XLTS n3047 n2769 n2849 gnd vdd NOR2XLTS
x462NOR2XLTS n3501 n3504 n3505 gnd vdd NOR2XLTS
x463NOR2XLTS n3505 n3506 n2753 gnd vdd NOR2XLTS
x464NOR2XLTS n3506 n2878 n2744 gnd vdd NOR2XLTS
x465NOR2XLTS n3504 n3507 n2724 gnd vdd NOR2XLTS
x466NOR2XLTS n3507 n2883 n2725 gnd vdd NOR2XLTS
x467NOR2XLTS n3224 n3225 n2715 gnd vdd NOR2XLTS
x468NOR2XLTS n3225 n2809 n2934 gnd vdd NOR2XLTS
x469NOR2XLTS n3223 n2813 n3167 gnd vdd NOR2XLTS
x470NOR2XLTS n3031 n3226 n3227 gnd vdd NOR2XLTS
x471NOR2XLTS n3228 n3230 n3231 gnd vdd NOR2XLTS
x472NOR2XLTS n3088 n2881 n2860 gnd vdd NOR2XLTS
x473NOR2XLTS n3230 n3235 n2796 gnd vdd NOR2XLTS
x474NOR2XLTS n3235 n2879 n2747 gnd vdd NOR2XLTS
x475NOR2XLTS n3237 n3238 n3239 gnd vdd NOR2XLTS
x476AND2XLTS n3244 n3245 n3242 gnd vdd AND2XLTS
x477INVXLTS n3004 n2839 gnd vdd INVXLTS
x478NOR2XLTS n3236 n3123 n3246 gnd vdd NOR2XLTS
x479NOR2XLTS n3246 n3109 n2734 gnd vdd NOR2XLTS
x480NOR2XLTS n3123 n3202 n2828 gnd vdd NOR2XLTS
x481NOR2XLTS n3248 n3438 n3439 gnd vdd NOR2XLTS
x482OR2XLTS n3440 n3441 n3439 gnd vdd OR2XLTS
x483NOR2XLTS n3449 n3450 n3451 gnd vdd NOR2XLTS
x484NOR2XLTS n3451 n3222 n2733 gnd vdd NOR2XLTS
x485NOR2XLTS n3450 n3171 n2793 gnd vdd NOR2XLTS
x486NOR2XLTS n3448 n3452 n3453 gnd vdd NOR2XLTS
x487NOR2XLTS n3454 n3456 n3457 gnd vdd NOR2XLTS
x488NOR2XLTS n3457 n2796 n2835 gnd vdd NOR2XLTS
x489NOR2XLTS n3456 n2767 n2814 gnd vdd NOR2XLTS
x490NOR2XLTS n3452 n2941 n2824 gnd vdd NOR2XLTS
x491NOR2XLTS n2941 n2852 n2855 gnd vdd NOR2XLTS
x492NOR2XLTS n3250 n3251 n3252 gnd vdd NOR2XLTS
x493NOR2XLTS n3249 n3259 n3260 gnd vdd NOR2XLTS
x494NOR2XLTS n3539 n3059 n3540 gnd vdd NOR2XLTS
x495NOR2XLTS n3541 n3545 n3546 gnd vdd NOR2XLTS
x496INVXLTS n3040 n3134 gnd vdd INVXLTS
x497NOR2XLTS n3544 n2873 n2779 gnd vdd NOR2XLTS
x498NOR2XLTS n3557 n3564 n3565 gnd vdd NOR2XLTS
x499NOR2XLTS n3564 n3572 n2757 gnd vdd NOR2XLTS
x500NOR2XLTS n3572 n2810 n3574 gnd vdd NOR2XLTS
x501NOR2XLTS n3538 n3058 n3575 gnd vdd NOR2XLTS
x502NOR2XLTS n3581 n3411 n3582 gnd vdd NOR2XLTS
x503NOR2XLTS n3582 n2822 n2771 gnd vdd NOR2XLTS
x504NOR2XLTS n3580 n3584 n3585 gnd vdd NOR2XLTS
x505NOR2XLTS n3585 n3171 n2805 gnd vdd NOR2XLTS
x506NOR2XLTS n3171 n2858 n2745 gnd vdd NOR2XLTS
x507NOR2XLTS n3584 n3588 n2720 gnd vdd NOR2XLTS
x508NOR2XLTS n3588 n2817 n2854 gnd vdd NOR2XLTS
x509NOR2XLTS n3269 n3270 n3271 gnd vdd NOR2XLTS
x510NOR2XLTS n3273 n2957 n2968 gnd vdd NOR2XLTS
x511NOR2XLTS n3275 n3276 n3277 gnd vdd NOR2XLTS
x512NOR2XLTS n3280 n3282 n3036 gnd vdd NOR2XLTS
x513NOR2XLTS n3036 n2800 n2814 gnd vdd NOR2XLTS
x514NOR2XLTS n3282 n2826 n2742 gnd vdd NOR2XLTS
x515NOR2XLTS n3274 n3283 n3284 gnd vdd NOR2XLTS
x516INVXLTS n3104 n3288 gnd vdd INVXLTS
x517NOR2XLTS n3132 n2912 n3289 gnd vdd NOR2XLTS
x518NOR2XLTS n3290 n3293 n3294 gnd vdd NOR2XLTS
x519NOR2XLTS n3294 n3109 n2766 gnd vdd NOR2XLTS
x520NOR2XLTS n3109 n2717 n2738 gnd vdd NOR2XLTS
x521NOR2XLTS n3293 n3295 n2861 gnd vdd NOR2XLTS
x522NOR2XLTS n3297 n3298 n3299 gnd vdd NOR2XLTS
x523NOR2XLTS n3299 n2954 n2831 gnd vdd NOR2XLTS
x524NOR2XLTS n3298 n2806 n2822 gnd vdd NOR2XLTS
x525NOR2XLTS n3296 n3300 n3301 gnd vdd NOR2XLTS
x526NOR2XLTS n3300 n2794 n2710 gnd vdd NOR2XLTS
x527NOR2XLTS n3272 n3305 n3306 gnd vdd NOR2XLTS
x528NOR2XLTS n3308 n3309 n3310 gnd vdd NOR2XLTS
x529NOR2XLTS n3310 n2716 n2805 gnd vdd NOR2XLTS
x530NOR2XLTS n3309 n2710 n2827 gnd vdd NOR2XLTS
x531NOR2XLTS n3307 n3311 n3312 gnd vdd NOR2XLTS
x532NOR2XLTS n3312 n2720 n2815 gnd vdd NOR2XLTS
x533NOR2XLTS n3311 n3151 n2775 gnd vdd NOR2XLTS
x534NOR2XLTS n3151 n2730 n3085 gnd vdd NOR2XLTS
x535NOR2XLTS n3314 n3315 n3316 gnd vdd NOR2XLTS
x536NOR2XLTS n3316 n3014 n2833 gnd vdd NOR2XLTS
x537NOR2XLTS n3014 n2693 n2765 gnd vdd NOR2XLTS
x538NOR2XLTS n3315 n3317 n2790 gnd vdd NOR2XLTS
x539NOR2XLTS n3317 n2701 n3257 gnd vdd NOR2XLTS
x540NOR2XLTS n3313 n3318 n3319 gnd vdd NOR2XLTS
x541NOR2XLTS n3319 n3320 n2727 gnd vdd NOR2XLTS
x542NOR2XLTS n3320 n2844 n2851 gnd vdd NOR2XLTS
x543NOR2XLTS n3318 n3321 n2800 gnd vdd NOR2XLTS
x544NOR2XLTS n3321 n2783 n2809 gnd vdd NOR2XLTS
x545OR2XLTS n3019 n3322 n3270 gnd vdd OR2XLTS
x546NOR2XLTS n3323 n3324 n3325 gnd vdd NOR2XLTS
x547NOR2XLTS n3325 n2762 n2742 gnd vdd NOR2XLTS
x548NOR2XLTS n3324 n2820 n2759 gnd vdd NOR2XLTS
x549NOR2XLTS n2960 n3326 n3327 gnd vdd NOR2XLTS
x550NOR2XLTS n2977 n2798 n2738 gnd vdd NOR2XLTS
x551NOR2XLTS n3331 n3334 n3335 gnd vdd NOR2XLTS
x552NOR2XLTS n3335 n3336 n2793 gnd vdd NOR2XLTS
x553NOR2XLTS n3336 n2882 n2870 gnd vdd NOR2XLTS
x554NOR2XLTS n3334 n3337 n2834 gnd vdd NOR2XLTS
x555NOR2XLTS n3337 n2718 n2816 gnd vdd NOR2XLTS
x556NOR2XLTS n3339 n3340 n3341 gnd vdd NOR2XLTS
x557INVXLTS n3023 n2740 gnd vdd INVXLTS
x558NOR2XLTS n3338 n3345 n3346 gnd vdd NOR2XLTS
x559NOR2XLTS n3350 n2871 n2859 gnd vdd NOR2XLTS
x560NOR2XLTS n3169 n2695 n2713 gnd vdd NOR2XLTS
x561INVXLTS n3097 n2792 gnd vdd INVXLTS
x562INVXLTS n2924 n2795 gnd vdd INVXLTS
x563NOR2XLTS n3295 n2797 n2842 gnd vdd NOR2XLTS
x564NOR2XLTS n2986 n3523 n3289 gnd vdd NOR2XLTS
x565NOR2XLTS n3222 n2811 n2714 gnd vdd NOR2XLTS
x566NOR2XLTS n2928 n3568 n3573 gnd vdd NOR2XLTS
x567NOR2XLTS n3357 n3363 n2788 gnd vdd NOR2XLTS
x568NOR2XLTS n3363 n2869 n2696 gnd vdd NOR2XLTS
x569INVXLTS n3006 n2824 gnd vdd INVXLTS
x570NOR2XLTS n3017 n3364 n3365 gnd vdd NOR2XLTS
x571NOR2XLTS n3366 n3368 n3369 gnd vdd NOR2XLTS
x572NOR2XLTS n3369 n2830 n2710 gnd vdd NOR2XLTS
x573NOR2XLTS n3368 n2803 n3167 gnd vdd NOR2XLTS
x574NOR2XLTS n3364 n2821 n2823 gnd vdd NOR2XLTS
x575NOR2XLTS n2955 n3371 n3372 gnd vdd NOR2XLTS
x576NOR2XLTS n3374 n3375 n3376 gnd vdd NOR2XLTS
x577NOR2XLTS n3376 n2835 n2731 gnd vdd NOR2XLTS
x578NOR2XLTS n3375 n2739 n2752 gnd vdd NOR2XLTS
x579NOR2XLTS n3373 n3377 n3378 gnd vdd NOR2XLTS
x580NOR2XLTS n3377 n2733 n2789 gnd vdd NOR2XLTS
x581NOR2XLTS n3381 n3382 n3383 gnd vdd NOR2XLTS
x582NOR2XLTS n3383 n2711 n2762 gnd vdd NOR2XLTS
x583NOR2XLTS n3382 n3384 n2791 gnd vdd NOR2XLTS
x584NOR2XLTS n3384 n2886 n2862 gnd vdd NOR2XLTS
x585NOR2XLTS n3380 n3385 n3386 gnd vdd NOR2XLTS
x586NOR2XLTS n3385 n3390 n2820 gnd vdd NOR2XLTS
x587NOR2XLTS n3390 n2729 n3115 gnd vdd NOR2XLTS
x588NOR2XLTS n3018 n3392 n3393 gnd vdd NOR2XLTS
x589NOR2XLTS n3561 n2909 n2912 gnd vdd NOR2XLTS
x590INVXLTS n3085 n2734 gnd vdd INVXLTS
x591NOR2XLTS n3399 n3402 n3403 gnd vdd NOR2XLTS
x592NOR2XLTS n3403 n3404 n2761 gnd vdd NOR2XLTS
x593NOR2XLTS n3402 n3405 n2728 gnd vdd NOR2XLTS
x594NOR2XLTS n3405 n2841 n2737 gnd vdd NOR2XLTS
x595NOR2XLTS n2965 n3406 n3407 gnd vdd NOR2XLTS
x596NOR2XLTS n3409 n3410 n3411 gnd vdd NOR2XLTS
x597NOR2XLTS n3411 n2802 n2834 gnd vdd NOR2XLTS
x598NOR2XLTS n3410 n2723 n2733 gnd vdd NOR2XLTS
x599NOR2XLTS n3408 n3412 n3413 gnd vdd NOR2XLTS
x600NOR2XLTS n3413 n2731 n2823 gnd vdd NOR2XLTS
x601INVXLTS n3304 n3398 gnd vdd INVXLTS
x602NOR2XLTS n3412 n2727 n2814 gnd vdd NOR2XLTS
x603NOR2XLTS n3415 n3416 n3417 gnd vdd NOR2XLTS
x604NOR2XLTS n3417 n3418 n2772 gnd vdd NOR2XLTS
x605NOR2XLTS n3051 n3461 n3583 gnd vdd NOR2XLTS
x606INVXLTS n3461 n3499 gnd vdd INVXLTS
x607NOR2XLTS n3418 n2857 n3288 gnd vdd NOR2XLTS
x608NOR2XLTS n2975 n3523 n3524 gnd vdd NOR2XLTS
x609NOR2XLTS n2939 n3556 n3289 gnd vdd NOR2XLTS
x610NOR2XLTS n3416 n3419 n2806 gnd vdd NOR2XLTS
x611NOR2XLTS n2946 n2903 n3398 gnd vdd NOR2XLTS
x612NOR2XLTS n3419 n2874 n2862 gnd vdd NOR2XLTS
x613NOR2XLTS n2933 n3526 n3527 gnd vdd NOR2XLTS
x614NOR2XLTS n2994 n3523 n3563 gnd vdd NOR2XLTS
x615OR2XLTS n2891 n2908 n3563 gnd vdd OR2XLTS
x616INVXLTS n3523 n3466 gnd vdd INVXLTS
x617NOR2XLTS n3414 n3420 n3421 gnd vdd NOR2XLTS
x618NOR2XLTS n2925 n3556 n3524 gnd vdd NOR2XLTS
x619NOR2XLTS n3077 n3526 n3556 gnd vdd NOR2XLTS
x620INVXLTS n3015 n2729 gnd vdd INVXLTS
x621NOR2XLTS n3161 n2708 n3583 gnd vdd NOR2XLTS
x622INVXLTS n3583 n3586 gnd vdd INVXLTS
x623NOR2XLTS n3586 n2893 n2906 gnd vdd NOR2XLTS
x624NOR2XLTS n3420 n3426 n3427 gnd vdd NOR2XLTS
x625AND2XLTS n2899 n2902 n3428 gnd vdd AND2XLTS
x626NOR2XLTS n3587 n2911 n3570 gnd vdd NOR2XLTS
x627INVXLTS n3560 n3568 gnd vdd INVXLTS
x628OR2XLTS n2896 n2891 n3568 gnd vdd OR2XLTS
x629NOR2XLTS n3446 n2896 n3289 gnd vdd NOR2XLTS
x630INVXLTS n3570 n2908 gnd vdd INVXLTS
x631NOR2XLTS n2935 n3526 n3578 gnd vdd NOR2XLTS
x632INVXLTS n3562 n2911 gnd vdd INVXLTS
x633INVXLTS n3526 n3370 gnd vdd INVXLTS
x634AND2XLTS n2890 n2909 n3370 gnd vdd AND2XLTS
x635NOR2XLTS n3003 n3004 n2875 gnd vdd NOR2XLTS
x636NOR2XLTS n3404 n2866 n2883 gnd vdd NOR2XLTS
x637NAND2X1TS n3131 n3499 n3500 gnd vdd NAND2X1TS
x638NOR2BX1TS n3500 n2906 n2894 gnd vdd NOR2BX1TS
x639NOR2X1TS n3499 n2902 n2900 gnd vdd NOR2X1TS
x640NOR2BX1TS n3466 n2897 n2913 gnd vdd NOR2BX1TS
x641NOR2BX1TS n3459 n2894 n2905 gnd vdd NOR2BX1TS
x642NOR2BX1TS n3555 n2900 n2902 gnd vdd NOR2BX1TS
x643NAND2X1TS n3556 n2912 n2896 gnd vdd NAND2X1TS
x644NOR2BX1TS n3460 n2903 n2899 gnd vdd NOR2BX1TS
x645NAND2X1TS n3289 n2890 n3570 gnd vdd NAND2X1TS
x646NAND2X1TS n3465 n3466 n2889 gnd vdd NAND2X1TS
x647NAND2X1TS d6 n2961 n2962 gnd vdd NAND2X1TS
x648NAND2X1TS n2964 n2965 n2966 gnd vdd NAND2X1TS
x649NAND2X1TS n2967 n2969 n2970 gnd vdd NAND2X1TS
x650NAND2X1TS n2972 n2973 n2974 gnd vdd NAND2X1TS
x651NAND2X1TS n2974 n2870 n2738 gnd vdd NAND2X1TS
x652NAND2X1TS n2973 n2817 n2976 gnd vdd NAND2X1TS
x653NAND2X1TS n2979 n2980 n2981 gnd vdd NAND2X1TS
x654NAND2BX1TS n2981 n2982 n2810 gnd vdd NAND2BX1TS
x655NAND2X1TS n2980 n2786 n2983 gnd vdd NAND2X1TS
x656NAND2X1TS n2983 n2780 n2758 gnd vdd NAND2X1TS
x657NAND2X1TS n2978 n2984 n2985 gnd vdd NAND2X1TS
x658NAND2X1TS n2985 n2859 n2987 gnd vdd NAND2X1TS
x659NAND2X1TS n2987 n2791 n2753 gnd vdd NAND2X1TS
x660NAND2X1TS n2984 n2844 n2989 gnd vdd NAND2X1TS
x661NAND2X1TS n2989 n2990 n2823 gnd vdd NAND2X1TS
x662NAND2X1TS n2991 n2992 n2993 gnd vdd NAND2X1TS
x663NAND2X1TS n2993 n2718 n2883 gnd vdd NAND2X1TS
x664NAND2X1TS n2992 n2994 n2769 gnd vdd NAND2X1TS
x665NAND2X1TS d5 n3026 n3027 gnd vdd NAND2X1TS
x666NAND2X1TS n3029 n3030 n3031 gnd vdd NAND2X1TS
x667NAND2X1TS n3033 n3034 n3035 gnd vdd NAND2X1TS
x668NAND2X1TS n3032 n3041 n3042 gnd vdd NAND2X1TS
x669NAND2X1TS n2976 n2727 n3045 gnd vdd NAND2X1TS
x670NAND2X1TS n3045 n2908 n3046 gnd vdd NAND2X1TS
x671NAND2X1TS n3467 n3468 n3469 gnd vdd NAND2X1TS
x672NAND2X1TS n3471 n3472 n3473 gnd vdd NAND2X1TS
x673NAND2X1TS n3473 n2873 n2751 gnd vdd NAND2X1TS
x674NAND2X1TS n3472 n2852 n3424 gnd vdd NAND2X1TS
x675NAND2X1TS n3475 n3476 n3477 gnd vdd NAND2X1TS
x676NAND2X1TS n3477 n3051 n3156 gnd vdd NAND2X1TS
x677NAND2X1TS n3476 n2810 n3478 gnd vdd NAND2X1TS
x678NAND2X1TS n3478 n2834 n2768 gnd vdd NAND2X1TS
x679NAND2X1TS n3474 n3479 n3480 gnd vdd NAND2X1TS
x680NAND2X1TS n3480 n2870 n3481 gnd vdd NAND2X1TS
x681NAND2X1TS n3481 n2827 n3482 gnd vdd NAND2X1TS
x682NAND2X1TS n3482 n2906 n2709 gnd vdd NAND2X1TS
x683NAND2X1TS n3052 n3054 n3055 gnd vdd NAND2X1TS
x684NAND2X1TS d4 n3060 n3061 gnd vdd NAND2X1TS
x685NAND2X1TS n3062 n3063 n3064 gnd vdd NAND2X1TS
x686NOR2BX1TS n3064 n2951 n3065 gnd vdd NOR2BX1TS
x687NAND2X1TS n3065 n2959 n3066 gnd vdd NAND2X1TS
x688NAND2X1TS n3068 n3069 n3070 gnd vdd NAND2X1TS
x689NAND2X1TS n3069 n2845 n2859 gnd vdd NAND2X1TS
x690NAND2X1TS n3099 n3100 n3101 gnd vdd NAND2X1TS
x691NAND2X1TS n3101 n2747 n3102 gnd vdd NAND2X1TS
x692NAND2X1TS n3102 n2760 n2826 gnd vdd NAND2X1TS
x693NAND2X1TS n3100 n2754 n3103 gnd vdd NAND2X1TS
x694NAND2X1TS n3103 n3104 n2758 gnd vdd NAND2X1TS
x695NAND2X1TS n3098 n3105 n3106 gnd vdd NAND2X1TS
x696NAND2X1TS n3112 n3113 n3114 gnd vdd NAND2X1TS
x697NAND2X1TS n3114 n2726 n2786 gnd vdd NAND2X1TS
x698NAND2X1TS n3113 n2769 n3115 gnd vdd NAND2X1TS
x699NAND2X1TS n3116 n3117 n3118 gnd vdd NAND2X1TS
x700NAND2X1TS n3120 n3121 n3122 gnd vdd NAND2X1TS
x701NAND2X1TS n3127 n3128 n3129 gnd vdd NAND2X1TS
x702NAND2X1TS n3129 n2871 n3130 gnd vdd NAND2X1TS
x703NAND2X1TS n3130 n2821 n2724 gnd vdd NAND2X1TS
x704NAND2X1TS n3128 n2770 n3132 gnd vdd NAND2X1TS
x705NAND2X1TS n3138 n3139 n3140 gnd vdd NAND2X1TS
x706NAND2X1TS n3140 n2862 n2852 gnd vdd NAND2X1TS
x707NAND2X1TS n3139 n2748 n2785 gnd vdd NAND2X1TS
x708NAND2X1TS n3137 n3142 n3143 gnd vdd NAND2X1TS
x709NAND2X1TS n3143 n2755 n2779 gnd vdd NAND2X1TS
x710NAND2X1TS n3142 n2865 n2848 gnd vdd NAND2X1TS
x711NAND2X1TS d7 n2914 n2915 gnd vdd NAND2X1TS
x712NAND2X1TS n2917 n2995 n2996 gnd vdd NAND2X1TS
x713NAND2X1TS n2998 n2999 n3000 gnd vdd NAND2X1TS
x714NAND2X1TS n3008 n3009 n3010 gnd vdd NAND2X1TS
x715NAND2X1TS n3010 n2725 n2713 gnd vdd NAND2X1TS
x716NAND2X1TS n2997 n3017 n3018 gnd vdd NAND2X1TS
x717NAND2X1TS n3020 n3021 n3022 gnd vdd NAND2X1TS
x718NAND2X1TS n3022 n2750 n2755 gnd vdd NAND2X1TS
x719NAND2X1TS n2916 n2918 n2919 gnd vdd NAND2X1TS
x720NAND2X1TS n2921 n2922 n2923 gnd vdd NAND2X1TS
x721NAND2X1TS n2923 n2729 n2817 gnd vdd NAND2X1TS
x722NAND2X1TS n2922 n2882 n2797 gnd vdd NAND2X1TS
x723NAND2X1TS n2920 n2926 n2927 gnd vdd NAND2X1TS
x724NAND2X1TS n2927 n2770 n2878 gnd vdd NAND2X1TS
x725NAND2X1TS n2926 n2811 n2702 gnd vdd NAND2X1TS
x726NAND2X1TS n2930 n2931 n2932 gnd vdd NAND2X1TS
x727NAND2X1TS n2932 n2863 n2934 gnd vdd NAND2X1TS
x728NAND2X1TS n2931 n2887 n2936 gnd vdd NAND2X1TS
x729NAND2X1TS n2929 n2937 n2938 gnd vdd NAND2X1TS
x730NAND2X1TS n2938 n2857 n2940 gnd vdd NAND2X1TS
x731NAND2X1TS n2940 n2941 n2791 gnd vdd NAND2X1TS
x732NAND2X1TS n2947 n2706 n2898 gnd vdd NAND2X1TS
x733NAND2X1TS n2949 n2950 n2951 gnd vdd NAND2X1TS
x734NAND2X1TS n3082 n3083 n3084 gnd vdd NAND2X1TS
x735NAND2X1TS n3084 n2816 n2778 gnd vdd NAND2X1TS
x736NAND2X1TS n3081 n3090 n3091 gnd vdd NAND2X1TS
x737NAND2X1TS n3091 n2845 n3092 gnd vdd NAND2X1TS
x738NAND2X1TS n3092 n2712 n2720 gnd vdd NAND2X1TS
x739NAND2X1TS n2953 n3144 n3145 gnd vdd NAND2X1TS
x740NAND2X1TS n3147 n3148 n3149 gnd vdd NAND2X1TS
x741NAND2X1TS n3149 n2875 n3150 gnd vdd NAND2X1TS
x742NAND2X1TS n3148 n2811 n2745 gnd vdd NAND2X1TS
x743NAND2X1TS n3153 n3154 n3155 gnd vdd NAND2X1TS
x744NAND2X1TS n3155 n2784 n3156 gnd vdd NAND2X1TS
x745NAND2X1TS n3156 n2954 n2781 gnd vdd NAND2X1TS
x746NAND2X1TS n3154 n2787 n3157 gnd vdd NAND2X1TS
x747NAND2X1TS n3157 n3158 n2727 gnd vdd NAND2X1TS
x748NAND2X1TS n3152 n3159 n3160 gnd vdd NAND2X1TS
x749NAND2X1TS n3160 n2855 n3162 gnd vdd NAND2X1TS
x750NAND2X1TS n3162 n2982 n2721 gnd vdd NAND2X1TS
x751NAND2X1TS n3159 n2879 n3163 gnd vdd NAND2X1TS
x752NAND2X1TS n3163 n2796 n2789 gnd vdd NAND2X1TS
x753NAND2X1TS n2948 n2955 n2956 gnd vdd NAND2X1TS
x754NAND2X1TS n2958 n2959 n2960 gnd vdd NAND2X1TS
x755NAND2X1TS n3072 n3073 n3074 gnd vdd NAND2X1TS
x756NAND2X1TS n3074 n2885 n2849 gnd vdd NAND2X1TS
x757NAND2X1TS n3073 n2798 n2725 gnd vdd NAND2X1TS
x758NAND2X1TS n3071 n3075 n3076 gnd vdd NAND2X1TS
x759NAND2X1TS n3076 n2865 n2842 gnd vdd NAND2X1TS
x760NAND2X1TS n3509 n3510 n3511 gnd vdd NAND2X1TS
x761NAND2X1TS n3513 n3514 n3515 gnd vdd NAND2X1TS
x762NAND2X1TS n3515 n2855 n3257 gnd vdd NAND2X1TS
x763NAND2X1TS n3520 n3521 n3522 gnd vdd NAND2X1TS
x764NAND2X1TS n3522 n2816 n2874 gnd vdd NAND2X1TS
x765NAND2X1TS n3521 n2869 n3458 gnd vdd NAND2X1TS
x766NAND2X1TS n3057 n3528 n3529 gnd vdd NAND2X1TS
x767NAND2X1TS n3534 n3535 n3342 gnd vdd NAND2X1TS
x768NAND2X1TS n3136 n2766 n2822 gnd vdd NAND2X1TS
x769NAND2X1TS n3168 n3169 n2788 gnd vdd NAND2X1TS
x770NAND2X1TS n3170 n2753 n2736 gnd vdd NAND2X1TS
x771NAND2X1TS n3070 n2717 n2887 gnd vdd NAND2X1TS
x772NAND2X1TS n3028 n3173 n3174 gnd vdd NAND2X1TS
x773NAND2X1TS n3176 n3430 n3431 gnd vdd NAND2X1TS
x774NAND2X1TS n3431 n2747 n2713 gnd vdd NAND2X1TS
x775NAND2X1TS n3433 n3434 n3435 gnd vdd NAND2X1TS
x776NAND2X1TS n3435 n2863 n2787 gnd vdd NAND2X1TS
x777NAND2X1TS n3434 n2797 n2860 gnd vdd NAND2X1TS
x778NAND2X1TS n3432 n3436 n3437 gnd vdd NAND2X1TS
x779NAND2X1TS n3437 n2924 n2866 gnd vdd NAND2X1TS
x780NAND2X1TS n3436 n2754 n2882 gnd vdd NAND2X1TS
x781NAND2X1TS n3175 n3177 n3178 gnd vdd NAND2X1TS
x782NAND2X1TS n3180 n3181 n3182 gnd vdd NAND2X1TS
x783NAND2X1TS n3182 n2885 n3183 gnd vdd NAND2X1TS
x784NAND2X1TS n3190 n3191 n3192 gnd vdd NAND2X1TS
x785NAND2X1TS n3192 n2939 n3193 gnd vdd NAND2X1TS
x786NAND2X1TS n3193 n2795 n2803 gnd vdd NAND2X1TS
x787NAND2X1TS n3191 n2867 n3194 gnd vdd NAND2X1TS
x788NAND2X1TS n3194 n2820 n2775 gnd vdd NAND2X1TS
x789NAND2X1TS n3197 n3198 n3199 gnd vdd NAND2X1TS
x790NAND2X1TS n3199 n2849 n2870 gnd vdd NAND2X1TS
x791NAND2X1TS n3179 n3204 n3205 gnd vdd NAND2X1TS
x792NAND2X1TS n3196 n3209 n3210 gnd vdd NAND2X1TS
x793NAND2X1TS n3166 n2800 n2743 gnd vdd NAND2X1TS
x794NAND2X1TS n3215 n3216 n3217 gnd vdd NAND2X1TS
x795NAND2BX1TS n3217 n2941 n2860 gnd vdd NAND2BX1TS
x796NAND2X1TS n3216 n2854 n3115 gnd vdd NAND2X1TS
x797NAND2X1TS n3203 n3487 n3488 gnd vdd NAND2X1TS
x798NAND2X1TS n3489 n3490 n3491 gnd vdd NAND2X1TS
x799NAND2X1TS n3491 n2817 n2886 gnd vdd NAND2X1TS
x800NAND2X1TS n3495 n3496 n3497 gnd vdd NAND2X1TS
x801NAND2X1TS n3497 n3004 n3150 gnd vdd NAND2X1TS
x802NAND2X1TS n3150 n3498 n2804 gnd vdd NAND2X1TS
x803NAND2BX1TS n3496 n3384 n2852 gnd vdd NAND2BX1TS
x804NAND2X1TS n3494 n3501 n3502 gnd vdd NAND2X1TS
x805NAND2X1TS n3502 n2730 n3503 gnd vdd NAND2X1TS
x806NAND2X1TS n3503 n3047 n2771 gnd vdd NAND2X1TS
x807NAND2X1TS n3220 n2885 n2783 gnd vdd NAND2X1TS
x808NAND2X1TS n3219 n2755 n2879 gnd vdd NAND2X1TS
x809NAND2X1TS n3221 n3109 n3222 gnd vdd NAND2X1TS
x810NAND2X1TS n2934 n2790 n2774 gnd vdd NAND2X1TS
x811NAND2X1TS n3227 n3228 n3229 gnd vdd NAND2X1TS
x812NAND2X1TS n3229 n3006 n2936 gnd vdd NAND2X1TS
x813NAND2X1TS n2936 n2988 n2731 gnd vdd NAND2X1TS
x814NAND2X1TS n3231 n3232 n3233 gnd vdd NAND2X1TS
x815NAND2BX1TS n3233 n3088 n2765 gnd vdd NAND2BX1TS
x816NAND2X1TS n3232 n2844 n3234 gnd vdd NAND2X1TS
x817NAND2X1TS n3234 n2782 n2716 gnd vdd NAND2X1TS
x818NAND2X1TS n3226 n3236 n3237 gnd vdd NAND2X1TS
x819NAND2X1TS n3239 n3240 n3241 gnd vdd NAND2X1TS
x820NAND2X1TS n3241 n2729 n2784 gnd vdd NAND2X1TS
x821NAND2X1TS n3238 n3242 n3243 gnd vdd NAND2X1TS
x822NAND2X1TS n3243 n2888 n2810 gnd vdd NAND2X1TS
x823NAND2X1TS n3245 n3004 n2770 gnd vdd NAND2X1TS
x824NAND2X1TS n3441 n3442 n3443 gnd vdd NAND2X1TS
x825NAND2X1TS n3443 n2883 n2737 gnd vdd NAND2X1TS
x826NAND2X1TS n3442 n2770 n3330 gnd vdd NAND2X1TS
x827NAND2X1TS n3440 n3444 n3445 gnd vdd NAND2X1TS
x828NAND2X1TS n3445 n3446 n2764 gnd vdd NAND2X1TS
x829NAND2X1TS n3444 n2862 n3447 gnd vdd NAND2X1TS
x830NAND2X1TS n3447 n2819 n2840 gnd vdd NAND2X1TS
x831NAND2X1TS n3438 n3448 n3449 gnd vdd NAND2X1TS
x832NAND2X1TS n3453 n3454 n3455 gnd vdd NAND2X1TS
x833NAND2X1TS n3455 n2887 n2785 gnd vdd NAND2X1TS
x834NAND2X1TS n3165 n3249 n3250 gnd vdd NAND2X1TS
x835NAND2X1TS n3252 n3253 n3254 gnd vdd NAND2X1TS
x836NAND2X1TS n3254 n2750 n2809 gnd vdd NAND2X1TS
x837NAND2X1TS n3253 n2875 n2714 gnd vdd NAND2X1TS
x838NAND2X1TS n3251 n3255 n3256 gnd vdd NAND2X1TS
x839NAND2X1TS n3256 n2754 n3257 gnd vdd NAND2X1TS
x840NAND2X1TS n3255 n2860 n3258 gnd vdd NAND2X1TS
x841NAND2X1TS n3260 n3261 n3262 gnd vdd NAND2X1TS
x842NAND2X1TS n3262 n2763 n3263 gnd vdd NAND2X1TS
x843NAND2X1TS n3263 n3040 n2782 gnd vdd NAND2X1TS
x844NAND2X1TS n3261 n3006 n3264 gnd vdd NAND2X1TS
x845NAND2X1TS n3264 n2792 n2776 gnd vdd NAND2X1TS
x846NAND2X1TS n3259 n3265 n3266 gnd vdd NAND2X1TS
x847NAND2X1TS n3266 n2751 n3267 gnd vdd NAND2X1TS
x848NAND2X1TS n3267 n2711 n2721 gnd vdd NAND2X1TS
x849NAND2X1TS n3265 n2886 n3268 gnd vdd NAND2X1TS
x850NAND2X1TS n3268 n2805 n2828 gnd vdd NAND2X1TS
x851NAND2X1TS n3247 n3538 n3539 gnd vdd NAND2X1TS
x852NAND2X1TS n3540 n3541 n3542 gnd vdd NAND2X1TS
x853NAND2X1TS n3542 n2756 n3543 gnd vdd NAND2X1TS
x854NAND2X1TS n3543 n3544 n2833 gnd vdd NAND2X1TS
x855NAND2X1TS n3546 n3547 n3548 gnd vdd NAND2X1TS
x856NAND2X1TS n3548 n2783 n3549 gnd vdd NAND2X1TS
x857NAND2X1TS n3549 n2739 n2767 gnd vdd NAND2X1TS
x858NAND2X1TS n3547 n2846 n3550 gnd vdd NAND2X1TS
x859NAND2X1TS n3550 n3040 n2733 gnd vdd NAND2X1TS
x860NAND2X1TS n3134 n2839 n2759 gnd vdd NAND2X1TS
x861NAND2X1TS n3545 n3551 n3552 gnd vdd NAND2X1TS
x862NAND2X1TS n3552 n2925 n3553 gnd vdd NAND2X1TS
x863NAND2X1TS n3553 n3169 n2775 gnd vdd NAND2X1TS
x864NAND2X1TS n3551 n2866 n3554 gnd vdd NAND2X1TS
x865NAND2X1TS n3554 n2732 n2827 gnd vdd NAND2X1TS
x866NAND2X1TS n3059 n3557 n3558 gnd vdd NAND2X1TS
x867NAND2X1TS n3558 n3097 n3559 gnd vdd NAND2X1TS
x868NAND2X1TS n3559 n3544 n2839 gnd vdd NAND2X1TS
x869NAND2X1TS n3565 n3566 n3567 gnd vdd NAND2X1TS
x870NAND2X1TS n3567 n2756 n3464 gnd vdd NAND2X1TS
x871NAND2X1TS n3464 n3015 n2766 gnd vdd NAND2X1TS
x872NAND2X1TS n3566 n3023 n3571 gnd vdd NAND2X1TS
x873NAND2X1TS n3571 n2803 n2752 gnd vdd NAND2X1TS
x874NAND2X1TS n3574 n2774 n2735 gnd vdd NAND2X1TS
x875NAND2X1TS n3575 n3576 n3577 gnd vdd NAND2X1TS
x876NAND2X1TS n3577 n2888 n2797 gnd vdd NAND2X1TS
x877NAND2X1TS n3576 n2858 n3579 gnd vdd NAND2X1TS
x878NAND2X1TS n3579 n2761 n2814 gnd vdd NAND2X1TS
x879NAND2X1TS n3058 n3580 n3581 gnd vdd NAND2X1TS
x880NAND2X1TS d1 n3060 n3269 gnd vdd NAND2X1TS
x881NAND2X1TS n3271 n3272 n3273 gnd vdd NAND2X1TS
x882NAND2X1TS n2968 n3274 n3275 gnd vdd NAND2X1TS
x883NAND2X1TS n3277 n3278 n3279 gnd vdd NAND2X1TS
x884NAND2X1TS n3279 n2867 n2798 gnd vdd NAND2X1TS
x885NAND2X1TS n3278 n2846 n2877 gnd vdd NAND2X1TS
x886NAND2X1TS n3276 n3280 n3281 gnd vdd NAND2X1TS
x887NAND2X1TS n3281 n2764 n2881 gnd vdd NAND2X1TS
x888NAND2X1TS n3284 n3285 n3286 gnd vdd NAND2X1TS
x889NAND2X1TS n3286 n2848 n3287 gnd vdd NAND2X1TS
x890NAND2X1TS n3287 n3104 n2739 gnd vdd NAND2X1TS
x891NAND2X1TS n3285 n3161 n3132 gnd vdd NAND2X1TS
x892NAND2X1TS n3283 n3290 n3291 gnd vdd NAND2X1TS
x893NAND2X1TS n3291 n2841 n3292 gnd vdd NAND2X1TS
x894NAND2X1TS n3292 n2837 n2823 gnd vdd NAND2X1TS
x895NAND2X1TS n2957 n3296 n3297 gnd vdd NAND2X1TS
x896NAND2X1TS n3301 n3302 n3303 gnd vdd NAND2X1TS
x897NAND2X1TS n3303 n3304 n2878 gnd vdd NAND2X1TS
x898NAND2X1TS n3302 n2765 n2986 gnd vdd NAND2X1TS
x899NAND2X1TS n3306 n3307 n3308 gnd vdd NAND2X1TS
x900NAND2X1TS n3305 n3313 n3314 gnd vdd NAND2X1TS
x901NAND2X1TS n3257 n2781 n2728 gnd vdd NAND2X1TS
x902NAND2X1TS n3322 n2960 n3323 gnd vdd NAND2X1TS
x903NAND2X1TS n3327 n3328 n3329 gnd vdd NAND2X1TS
x904NAND2X1TS n3329 n2701 n2737 gnd vdd NAND2X1TS
x905NAND2X1TS n3328 n2854 n3330 gnd vdd NAND2X1TS
x906NAND2X1TS n3326 n3331 n3332 gnd vdd NAND2X1TS
x907NAND2X1TS n3332 n2858 n3333 gnd vdd NAND2X1TS
x908NAND2X1TS n3333 n2977 n2830 gnd vdd NAND2X1TS
x909NAND2X1TS n3019 n3338 n3339 gnd vdd NAND2X1TS
x910NAND2X1TS n3341 n3240 n3342 gnd vdd NAND2X1TS
x911NAND2X1TS n3342 n2886 n2769 gnd vdd NAND2X1TS
x912NAND2X1TS n3240 n3023 n2786 gnd vdd NAND2X1TS
x913NAND2X1TS n3340 n3343 n3344 gnd vdd NAND2X1TS
x914NAND2X1TS n3344 n3097 n3330 gnd vdd NAND2X1TS
x915NAND2X1TS n3330 n2704 n2742 gnd vdd NAND2X1TS
x916NAND2X1TS n3343 n2857 n2763 gnd vdd NAND2X1TS
x917NAND2X1TS n3346 n3347 n3348 gnd vdd NAND2X1TS
x918NAND2X1TS n3348 n2809 n3349 gnd vdd NAND2X1TS
x919NAND2X1TS n3349 n3350 n2781 gnd vdd NAND2X1TS
x920NAND2X1TS n3347 n2877 n3351 gnd vdd NAND2X1TS
x921NAND2X1TS n3351 n3169 n2802 gnd vdd NAND2X1TS
x922NAND2X1TS n3345 n3352 n3353 gnd vdd NAND2X1TS
x923NAND2X1TS n3353 n2924 n3354 gnd vdd NAND2X1TS
x924NAND2X1TS n3354 n2838 n2767 gnd vdd NAND2X1TS
x925NAND2X1TS n3352 n2744 n3355 gnd vdd NAND2X1TS
x926NAND2X1TS n3355 n3295 n2831 gnd vdd NAND2X1TS
x927NAND2X1TS n3013 n2707 n3460 gnd vdd NAND2X1TS
x928NAND2X1TS n3356 n2820 n2792 gnd vdd NAND2X1TS
x929NAND2X1TS n3358 n3359 n3360 gnd vdd NAND2X1TS
x930NAND2X1TS n3360 n2798 n3361 gnd vdd NAND2X1TS
x931NAND2X1TS n3361 n2800 n2757 gnd vdd NAND2X1TS
x932NAND2X1TS n3573 n2911 n2908 gnd vdd NAND2X1TS
x933NAND2X1TS n3359 n2726 n3362 gnd vdd NAND2X1TS
x934NAND2X1TS n3362 n2829 n2735 gnd vdd NAND2X1TS
x935NAND2X1TS n3365 n3366 n3367 gnd vdd NAND2X1TS
x936NAND2X1TS n3367 n2844 n2865 gnd vdd NAND2X1TS
x937NAND2X1TS n3167 n3370 n2897 gnd vdd NAND2X1TS
x938NAND2X1TS n3372 n3373 n3374 gnd vdd NAND2X1TS
x939NAND2X1TS n2988 n3499 n2706 gnd vdd NAND2X1TS
x940NAND2X1TS n3378 n3379 n3244 gnd vdd NAND2X1TS
x941NAND2X1TS n3244 n2869 n2851 gnd vdd NAND2X1TS
x942NAND2X1TS n3379 n2881 n2848 gnd vdd NAND2X1TS
x943NAND2X1TS n3125 n3459 n2709 gnd vdd NAND2X1TS
x944NAND2X1TS n3371 n3380 n3381 gnd vdd NAND2X1TS
x945NAND2X1TS n3386 n3387 n3388 gnd vdd NAND2X1TS
x946NAND2X1TS n3388 n2866 n3389 gnd vdd NAND2X1TS
x947NAND2X1TS n3389 n2794 n2829 gnd vdd NAND2X1TS
x948NAND2X1TS n3089 n3459 n3428 gnd vdd NAND2X1TS
x949NAND2X1TS n3387 n2874 n3258 gnd vdd NAND2X1TS
x950NAND2X1TS n3258 n2795 n2723 gnd vdd NAND2X1TS
x951NAND2X1TS n3115 n2740 n2838 gnd vdd NAND2X1TS
x952NAND2X1TS n3391 n2730 n2845 gnd vdd NAND2X1TS
x953NAND2X1TS n3393 n3394 n3395 gnd vdd NAND2X1TS
x954NAND2X1TS n3395 n2714 n3396 gnd vdd NAND2X1TS
x955NAND2X1TS n3396 n2837 n2715 gnd vdd NAND2X1TS
x956NAND2X1TS n2954 n3560 n3561 gnd vdd NAND2X1TS
x957NAND2X1TS n3394 n2698 n3397 gnd vdd NAND2X1TS
x958NAND2X1TS n3397 n3398 n2772 gnd vdd NAND2X1TS
x959NAND2X1TS n3392 n3399 n3400 gnd vdd NAND2X1TS
x960NAND2X1TS n3400 n2725 n3401 gnd vdd NAND2X1TS
x961NAND2X1TS n3401 n2793 n2806 gnd vdd NAND2X1TS
x962NAND2X1TS n3407 n3408 n3409 gnd vdd NAND2X1TS
x963NAND2X1TS n3096 n2707 n3428 gnd vdd NAND2X1TS
x964NAND2X1TS n3406 n3414 n3415 gnd vdd NAND2X1TS
x965NAND2X1TS n3288 n2697 n2722 gnd vdd NAND2X1TS
x966NAND2X1TS n3398 n2899 n3586 gnd vdd NAND2X1TS
x967NAND2X1TS n3527 n2912 n2895 gnd vdd NAND2X1TS
x968NAND2X1TS n3421 n3422 n3423 gnd vdd NAND2X1TS
x969NAND2X1TS n3423 n2738 n3424 gnd vdd NAND2X1TS
x970NAND2X1TS n3424 n2801 n2719 gnd vdd NAND2X1TS
x971NAND2X1TS n3524 n2909 n2889 gnd vdd NAND2X1TS
x972NAND2X1TS n3080 n3555 n3459 gnd vdd NAND2X1TS
x973NAND2X1TS n3422 n2854 n3425 gnd vdd NAND2X1TS
x974NAND2X1TS n3425 n2801 n2780 gnd vdd NAND2X1TS
x975NAND2X1TS n3569 n2911 n3570 gnd vdd NAND2X1TS
x976NAND2X1TS n3427 n2893 n3428 gnd vdd NAND2X1TS
x977MXI2X1TS n3426 n3429 n2744 n2905 gnd vdd MXI2X1TS
x978NAND2X1TS n2945 n3560 n3587 gnd vdd NAND2X1TS
x979NAND2X1TS n3429 n2728 n2824 gnd vdd NAND2X1TS
x980NAND2X1TS n3578 n2895 n3562 gnd vdd NAND2X1TS
.ends
