library verilog;
use verilog.vl_types.all;
entity prechargeinput_tb is
end prechargeinput_tb;
