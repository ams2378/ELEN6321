.SUBCKT CLKBUFX2TS A Y VSS VDD
X0 VDD nmin Y VDD LPPFET W=1.3U L=0.12U M=1
X1 Y nmin VSS VSS LPNFET W=0.48U L=0.12U M=1
X2 VDD A nmin VDD LPPFET W=0.54U L=0.12U M=1
X3 nmin A VSS VSS LPNFET W=0.2U L=0.12U M=1
.ENDS CLKBUFX2TS

.SUBCKT INVXLTS A Y  VSS VDD
X0 VDD A Y VDD LPPFET W=0.34U L=0.12U M=1
X1 Y A VSS VSS LPNFET W=0.24U L=0.12U M=1
.ENDS INVXLTS

.SUBCKT DFFSXLTS CK D Q QN SN  VSS VDD
X0 net52 s VDD VDD LPPFET W=0.28U L=0.12U M=1
X1 m SN VDD VDD LPPFET W=0.28U L=0.12U M=1
X10 net82 c m VSS LPNFET W=0.2U L=0.12U M=1
X11 hnet21 D VSS VSS LPNFET W=0.2U L=0.12U M=1
X12 pm cn hnet21 VSS LPNFET W=0.2U L=0.12U M=1
X13 hnet23 c pm VDD LPPFET W=0.28U L=0.12U M=1
X14 VDD D hnet23 VDD LPPFET W=0.28U L=0.12U M=1
X15 hnet27 m VSS VSS LPNFET W=0.22U L=0.12U M=1
X16 pm c hnet27 VSS LPNFET W=0.22U L=0.12U M=1
X17 hnet29 cn pm VDD LPPFET W=0.28U L=0.12U M=1
X18 VDD m hnet29 VDD LPPFET W=0.28U L=0.12U M=1
X19 VDD s net91 VDD LPPFET W=0.28U L=0.12U M=1
X2 m pm VDD VDD LPPFET W=0.28U L=0.12U M=1
X20 net91 s VSS VSS LPNFET W=0.2U L=0.12U M=1
X21 VDD s Q VDD LPPFET W=0.34U L=0.12U M=1
X22 Q s VSS VSS LPNFET W=0.24U L=0.12U M=1
X23 VDD net82 s VDD LPPFET W=0.28U L=0.12U M=1
X24 s net82 VSS VSS LPNFET W=0.2U L=0.12U M=1
X25 VDD net91 QN VDD LPPFET W=0.34U L=0.12U M=1
X26 QN net91 VSS VSS LPNFET W=0.24U L=0.12U M=1
X27 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1
X28 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1
X29 VDD CK cn VDD LPPFET W=0.42U L=0.12U M=1
X3 net82 SN VDD VDD LPPFET W=0.28U L=0.12U M=1
X30 cn CK VSS VSS LPNFET W=0.3U L=0.12U M=1
X4 net82 c net52 VDD LPPFET W=0.28U L=0.12U M=1
X5 net82 cn m VDD LPPFET W=0.28U L=0.12U M=1
X6 m pm net76 VSS LPNFET W=0.3U L=0.12U M=1
X7 net73 s net76 VSS LPNFET W=0.2U L=0.12U M=1
X8 net76 SN VSS VSS LPNFET W=0.4U L=0.12U M=1
X9 net82 cn net73 VSS LPNFET W=0.2U L=0.12U M=1
.ENDS DFFSXLTS

.SUBCKT XOR2X1TS A B Y VSS VDD
X0 Y A net35 VDD LPPFET W=0.76U L=0.12U M=1
X1 Y nmin1 nmin2 VDD LPPFET W=0.78U L=0.12U M=1
X2 Y nmin1 net35 VSS LPNFET W=0.56U L=0.12U M=1
X3 Y A nmin2 VSS LPNFET W=0.54U L=0.12U M=1
X4 VDD A nmin1 VDD LPPFET W=0.3U L=0.12U M=1
X5 nmin1 A VSS VSS LPNFET W=0.22U L=0.12U M=1
X6 VDD nmin2 net35 VDD LPPFET W=0.76U L=0.12U M=1
X7 net35 nmin2 VSS VSS LPNFET W=0.56U L=0.12U M=1
X8 VDD B nmin2 VDD LPPFET W=0.78U L=0.12U M=1
X9 nmin2 B VSS VSS LPNFET W=0.54U L=0.12U M=1
.ENDS XOR2X1TS
