*.GLOBAL VDD VSS VSS1 
*.SCALE METER 

**** 
*.SUBCKT ACCSHCINX2TS CO0 CO1 A B CI0N CI1N 
.SUBCKT ACCSHCINX2TS CO0 CO1 A B CI0N CI1N VSS VDD
X0 CO1 net124 net137 VDD LPPFET W=1.3U L=0.12U M=1 
X1 CO1 net118 nmcin1n VDD LPPFET W=1.3U L=0.12U M=1 
X10 CO0 net118 net125 VSS LPNFET W=0.92U L=0.12U M=1 
X11 CO0 net124 nmcin0n VSS LPNFET W=0.92U L=0.12U M=1 
X12 net118 B net135 VSS LPNFET W=0.9U L=0.12U M=1 
X13 net118 nmb nma VSS LPNFET W=0.84U L=0.12U M=1 
X14 net124 B nma VSS LPNFET W=0.86U L=0.12U M=1 
X15 net124 nmb net135 VSS LPNFET W=0.92U L=0.12U M=1 
X16 VDD nmb net125 VDD LPPFET W=1.3U L=0.12U M=1 
X17 net125 nmb VSS VSS LPNFET W=0.92U L=0.12U M=1 
X18 VDD CI1N nmcin1n VDD LPPFET W=1.3U L=0.12U M=1 
X19 nmcin1n CI1N VSS VSS LPNFET W=0.92U L=0.12U M=1
X2 CO0 net124 net125 VDD LPPFET W=1.3U L=0.12U M=1 
X20 VDD CI0N nmcin0n VDD LPPFET W=1.3U L=0.12U M=1 
X21 nmcin0n CI0N VSS VSS LPNFET W=0.92U L=0.12U M=1 
X22 VDD B nmb VDD LPPFET W=1.28U L=0.12U M=1 
X23 nmb B VSS VSS LPNFET W=0.92U L=0.12U M=1 
X24 VDD A nma VDD LPPFET W=1.3U L=0.12U M=1 
X25 nma A VSS VSS LPNFET W=0.9U L=0.12U M=1 
X26 VDD nma net135 VDD LPPFET W=1.24U L=0.12U M=1 
X27 net135 nma VSS VSS LPNFET W=0.9U L=0.12U M=1 
X28 VDD nma net137 VDD LPPFET W=1.24U L=0.12U M=1 
X29 net137 nma VSS VSS LPNFET W=0.9U L=0.12U M=1 
X3 CO0 net118 nmcin0n VDD LPPFET W=1.3U L=0.12U M=1 
X4 net118 nmb net135 VDD LPPFET W=1.24U L=0.12U M=1 
X5 net118 B nma VDD LPPFET W=1.28U L=0.12U M=1 
X6 net124 nmb nma VDD LPPFET W=1.28U L=0.12U M=1 
X7 net124 B net135 VDD LPPFET W=1.28U L=0.12U M=1 
X8 CO1 net118 net137 VSS LPNFET W=0.86U L=0.12U M=1 
X9 CO1 net124 nmcin1n VSS LPNFET W=0.86U L=0.12U M=1 
.ENDS ACCSHCINX2TS 

**** 
*.SUBCKT ACCSHCINX4TS CO0 CO1 A B CI0N CI1N 
.SUBCKT ACCSHCINX4TS CO0 CO1 A B CI0N CI1N VSS VDD
X0 CO1 net126 net139 VDD LPPFET W=1.2U L=0.12U M=1 
X1 CO1 net120 net129 VDD LPPFET W=2.6U L=0.12U M=1 
X10 CO0 net120 net127 VSS LPNFET W=0.92U L=0.12U M=1 
X11 CO0 net126 net131 VSS LPNFET W=1.84U L=0.12U M=1 
X12 net120 B net137 VSS LPNFET W=0.9U L=0.12U M=1 
X13 net120 net133 net140 VSS LPNFET W=0.84U L=0.12U M=1 
X14 net126 B net140 VSS LPNFET W=0.86U L=0.12U M=1 
X15 net126 net133 net137 VSS LPNFET W=0.92U L=0.12U M=1 
X16 VDD net133 net127 VDD LPPFET W=1.3U L=0.12U M=1 
X17 net127 net133 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X18 VDD CI1N net129 VDD LPPFET W=2.6U L=0.12U M=1 
X19 net129 CI1N VSS VSS LPNFET W=1.84U L=0.12U M=1 
X2 CO0 net126 net127 VDD LPPFET W=1.2U L=0.12U M=1 
X20 VDD CI0N net131 VDD LPPFET W=2.6U L=0.12U M=1 
X21 net131 CI0N VSS VSS LPNFET W=1.84U L=0.12U M=1 
X22 VDD B net133 VDD LPPFET W=1.28U L=0.12U M=1 
X23 net133 B VSS VSS LPNFET W=0.92U L=0.12U M=1 
X24 VDD A net140 VDD LPPFET W=1.3U L=0.12U M=1 
X25 net140 A VSS VSS LPNFET W=0.9U L=0.12U M=1 
X26 VDD net140 net137 VDD LPPFET W=1.24U L=0.12U M=1 
X27 net137 net140 VSS VSS LPNFET W=0.9U L=0.12U M=1 
X28 VDD net140 net139 VDD LPPFET W=1.24U L=0.12U M=1 
X29 net139 net140 VSS VSS LPNFET W=0.9U L=0.12U M=1 
X3 CO0 net120 net131 VDD LPPFET W=2.34U L=0.12U M=1 
X4 net120 net133 net137 VDD LPPFET W=1.24U L=0.12U M=1 
X5 net120 B net140 VDD LPPFET W=1.28U L=0.12U M=1 
X6 net126 net133 net140 VDD LPPFET W=1.28U L=0.12U M=1 
X7 net126 B net137 VDD LPPFET W=1.28U L=0.12U M=1 
X8 CO1 net120 net139 VSS LPNFET W=0.92U L=0.12U M=1 
X9 CO1 net126 net129 VSS LPNFET W=1.72U L=0.12U M=1 
.ENDS ACCSHCINX4TS 

**** 
*.SUBCKT ACCSHCONX2TS CO0N CO1N A B CI0 CI1 
.SUBCKT ACCSHCONX2TS CO0N CO1N A B CI0 CI1 VSS VDD
X0 CO1N net99 net97 VDD LPPFET W=1.3U L=0.12U M=1 
X1 CO1N net96 nmcin1 VDD LPPFET W=1.28U L=0.12U M=1 
X10 net96 B net109 VSS LPNFET W=0.86U L=0.12U M=1 
X11 net96 nmb nma VSS LPNFET W=0.92U L=0.12U M=1 
X12 VDD B net97 VDD LPPFET W=1.3U L=0.12U M=1 
X13 net97 B VSS VSS LPNFET W=0.88U L=0.12U M=1 
X14 VDD net96 net99 VDD LPPFET W=1.28U L=0.12U M=1 
X15 net99 net96 VSS VSS LPNFET W=0.9U L=0.12U M=1 
X16 VDD CI1 nmcin1 VDD LPPFET W=1.3U L=0.12U M=1 
X17 nmcin1 CI1 VSS VSS LPNFET W=0.86U L=0.12U M=1 
X18 VDD CI0 nmcin0 VDD LPPFET W=1.3U L=0.12U M=1 
X19 nmcin0 CI0 VSS VSS LPNFET W=0.86U L=0.12U M=1 
X2 CO0N net99 net111 VDD LPPFET W=1.28U L=0.12U M=1 
X20 VDD B nmb VDD LPPFET W=1.3U L=0.12U M=1 
X21 nmb B VSS VSS LPNFET W=0.88U L=0.12U M=1 
X22 VDD A nma VDD LPPFET W=1.3U L=0.12U M=1 
X23 nma A VSS VSS LPNFET W=0.86U L=0.12U M=1 
X24 VDD nma net109 VDD LPPFET W=1.3U L=0.12U M=1 
X25 net109 nma VSS VSS LPNFET W=0.86U L=0.12U M=1 
X26 VDD A net111 VDD LPPFET W=1.3U L=0.12U M=1 
X27 net111 A VSS VSS LPNFET W=0.92U L=0.12U M=1 
X3 CO0N net96 nmcin0 VDD LPPFET W=1.2U L=0.12U M=1 
X4 net96 nmb net109 VDD LPPFET W=1.3U L=0.12U M=1 
X5 net96 B nma VDD LPPFET W=1.3U L=0.12U M=1 
X6 CO1N net96 net97 VSS LPNFET W=0.92U L=0.12U M=1 
X7 CO1N net99 nmcin1 VSS LPNFET W=0.88U L=0.12U M=1 
X8 CO0N net96 net111 VSS LPNFET W=0.88U L=0.12U M=1 
X9 CO0N net99 nmcin0 VSS LPNFET W=0.86U L=0.12U M=1 
.ENDS ACCSHCONX2TS 

**** 
*.SUBCKT ACCSHCONX4TS CO0N CO1N A B CI0 CI1 
.SUBCKT ACCSHCONX4TS CO0N CO1N A B CI0 CI1 VSS VDD
X0 CO1N net99 net97 VDD LPPFET W=1.3U L=0.12U M=1 
X1 CO1N net96 nmcin1 VDD LPPFET W=2.5U L=0.12U M=1 
X10 net96 B net109 VSS LPNFET W=0.86U L=0.12U M=1 
X11 net96 nmb nma VSS LPNFET W=0.92U L=0.12U M=1 
X12 VDD B net97 VDD LPPFET W=1.3U L=0.12U M=1 
X13 net97 B VSS VSS LPNFET W=0.88U L=0.12U M=1 
X14 VDD net96 net99 VDD LPPFET W=1.24U L=0.12U M=1 
X15 net99 net96 VSS VSS LPNFET W=0.9U L=0.12U M=1 
X16 VDD CI1 nmcin1 VDD LPPFET W=2.6U L=0.12U M=1 
X17 nmcin1 CI1 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X18 VDD CI0 nmcin0 VDD LPPFET W=2.6U L=0.12U M=1 
X19 nmcin0 CI0 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X2 CO0N net99 net111 VDD LPPFET W=1.22U L=0.12U M=1 
X20 VDD B nmb VDD LPPFET W=1.3U L=0.12U M=1 
X21 nmb B VSS VSS LPNFET W=0.88U L=0.12U M=1 
X22 VDD A nma VDD LPPFET W=1.3U L=0.12U M=1 
X23 nma A VSS VSS LPNFET W=0.86U L=0.12U M=1 
X24 VDD nma net109 VDD LPPFET W=1.3U L=0.12U M=1 
X25 net109 nma VSS VSS LPNFET W=0.86U L=0.12U M=1 
X26 VDD A net111 VDD LPPFET W=1.3U L=0.12U M=1 
X27 net111 A VSS VSS LPNFET W=0.92U L=0.12U M=1 
X3 CO0N net96 nmcin0 VDD LPPFET W=2.5U L=0.12U M=1 
X4 net96 nmb net109 VDD LPPFET W=1.3U L=0.12U M=1 
X5 net96 B nma VDD LPPFET W=1.3U L=0.12U M=1 
X6 CO1N net96 net97 VSS LPNFET W=0.92U L=0.12U M=1 
X7 CO1N net99 nmcin1 VSS LPNFET W=1.82U L=0.12U M=1 
X8 CO0N net96 net111 VSS LPNFET W=0.88U L=0.12U M=1 
X9 CO0N net99 nmcin0 VSS LPNFET W=1.82U L=0.12U M=1 
.ENDS ACCSHCONX4TS 

**** 
*.SUBCKT ACCSIHCONX2TS CO0N CO1N A B 
.SUBCKT ACCSIHCONX2TS CO0N CO1N A B VSS VDD
X0 CO1N B VSS VSS LPNFET W=0.72U L=0.12U M=1 
X1 CO1N A VSS VSS LPNFET W=0.72U L=0.12U M=1 
X2 VDD B hnet8 VDD LPPFET W=1.3U L=0.12U M=1 
X3 hnet8 A CO1N VDD LPPFET W=1.3U L=0.12U M=1 
X4 hnet16 A VSS VSS LPNFET W=0.92U L=0.12U M=1 
X5 CO0N B hnet16 VSS LPNFET W=0.92U L=0.12U M=1 
X6 VDD A CO0N VDD LPPFET W=0.96U L=0.12U M=1 
X7 VDD B CO0N VDD LPPFET W=0.96U L=0.12U M=1 
.ENDS ACCSIHCONX2TS 

**** 
*.SUBCKT ACCSIHCONX4TS CO0N CO1N A B 
.SUBCKT ACCSIHCONX4TS CO0N CO1N A B VSS VDD
X0 CO1N B VSS VSS LPNFET W=1.32U L=0.12U M=1 
X1 CO1N A VSS VSS LPNFET W=1.32U L=0.12U M=1 
X10 VDD A CO0N VDD LPPFET W=1.88U L=0.12U M=1 
X11 VDD B CO0N VDD LPPFET W=1.88U L=0.12U M=1 
X2 VDD B hnet9 VDD LPPFET W=1.3U L=0.12U M=1 
X3 hnet9 A CO1N VDD LPPFET W=1.3U L=0.12U M=1 
X4 VDD B hnet7 VDD LPPFET W=1.3U L=0.12U M=1 
X5 hnet7 A CO1N VDD LPPFET W=1.3U L=0.12U M=1 
X6 hnet18 A VSS VSS LPNFET W=0.9U L=0.12U M=1 
X7 CO0N B hnet18 VSS LPNFET W=0.9U L=0.12U M=1 
X8 hnet14 A VSS VSS LPNFET W=0.9U L=0.12U M=1 
X9 CO0N B hnet14 VSS LPNFET W=0.9U L=0.12U M=1 
.ENDS ACCSIHCONX4TS 

**** 
*.SUBCKT ACHCINX2TS CO A B CIN 
.SUBCKT ACHCINX2TS CO A B CIN VSS VDD
X0 VDD nmb net59 VDD LPPFET W=1.3U L=0.12U M=1 
X1 net59 nmb VSS VSS LPNFET W=0.92U L=0.12U M=1 
X10 CO net104 net59 VDD LPPFET W=1.3U L=0.12U M=1 
X11 CO net98 nmcinn VDD LPPFET W=1.22U L=0.12U M=1 
X12 net98 nmb net67 VDD LPPFET W=1.02U L=0.12U M=1 
X13 net98 B nma VDD LPPFET W=1.3U L=0.12U M=1 
X14 net104 nmb nma VDD LPPFET W=1.16U L=0.12U M=1 
X15 net104 B net67 VDD LPPFET W=1.02U L=0.12U M=1 
X16 CO net98 net59 VSS LPNFET W=0.92U L=0.12U M=1 
X17 CO net104 nmcinn VSS LPNFET W=0.92U L=0.12U M=1 
X18 net98 B net67 VSS LPNFET W=0.74U L=0.12U M=1 
X19 net98 nmb nma VSS LPNFET W=0.84U L=0.12U M=1 
X2 VDD CIN nmcinn VDD LPPFET W=1.22U L=0.12U M=1 
X20 net104 B nma VSS LPNFET W=0.88U L=0.12U M=1 
X21 net104 nmb net67 VSS LPNFET W=0.76U L=0.12U M=1 
X3 nmcinn CIN VSS VSS LPNFET W=0.92U L=0.12U M=1 
X4 VDD B nmb VDD LPPFET W=1.3U L=0.12U M=1 
X5 nmb B VSS VSS LPNFET W=0.92U L=0.12U M=1 
X6 VDD A nma VDD LPPFET W=1.3U L=0.12U M=1 
X7 nma A VSS VSS LPNFET W=0.92U L=0.12U M=1 
X8 VDD nma net67 VDD LPPFET W=1.02U L=0.12U M=1 
X9 net67 nma VSS VSS LPNFET W=0.74U L=0.12U M=1 
.ENDS ACHCINX2TS 

**** 
*.SUBCKT ACHCINX4TS CO A B CIN 
.SUBCKT ACHCINX4TS CO A B CIN VSS VDD
X0 VDD net64 net60 VDD LPPFET W=1.3U L=0.12U M=1 
X1 net60 net64 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X10 CO net105 net60 VDD LPPFET W=1.3U L=0.12U M=1 
X11 CO net99 net62 VDD LPPFET W=2.36U L=0.12U M=1 
X12 net99 net64 net68 VDD LPPFET W=1.24U L=0.12U M=1 
X13 net99 B net66 VDD LPPFET W=1.3U L=0.12U M=1 
X14 net105 net64 net66 VDD LPPFET W=1.28U L=0.12U M=1 
X15 net105 B net68 VDD LPPFET W=1.28U L=0.12U M=1 
X16 CO net99 net60 VSS LPNFET W=0.92U L=0.12U M=1 
X17 CO net105 net62 VSS LPNFET W=1.84U L=0.12U M=1 
X18 net99 B net68 VSS LPNFET W=0.92U L=0.12U M=1 
X19 net99 net64 net66 VSS LPNFET W=0.88U L=0.12U M=1 
X2 VDD CIN net62 VDD LPPFET W=2.36U L=0.12U M=1 
X20 net105 B net66 VSS LPNFET W=0.86U L=0.12U M=1 
X21 net105 net64 net68 VSS LPNFET W=0.92U L=0.12U M=1 
X3 net62 CIN VSS VSS LPNFET W=1.84U L=0.12U M=1 
X4 VDD B net64 VDD LPPFET W=1.3U L=0.12U M=1 
X5 net64 B VSS VSS LPNFET W=0.92U L=0.12U M=1 
X6 VDD A net66 VDD LPPFET W=1.3U L=0.12U M=1 
X7 net66 A VSS VSS LPNFET W=0.92U L=0.12U M=1 
X8 VDD net66 net68 VDD LPPFET W=1.24U L=0.12U M=1 
X9 net68 net66 VSS VSS LPNFET W=0.92U L=0.12U M=1 
.ENDS ACHCINX4TS 

**** 
*.SUBCKT ACHCONX2TS CON A B CI 
.SUBCKT ACHCONX2TS CON A B CI VSS VDD
X0 VDD B nmb VDD LPPFET W=1.3U L=0.12U M=1 
X1 nmb B VSS VSS LPNFET W=0.92U L=0.12U M=1 
X10 CON net104 net63 VDD LPPFET W=1.3U L=0.12U M=1 
X11 CON net98 nmcin VDD LPPFET W=1.22U L=0.12U M=1 
X12 net98 nmb net67 VDD LPPFET W=1.02U L=0.12U M=1 
X13 net98 B nma VDD LPPFET W=1.3U L=0.12U M=1 
X14 net104 nmb nma VDD LPPFET W=1.16U L=0.12U M=1 
X15 net104 B net67 VDD LPPFET W=1.02U L=0.12U M=1 
X16 CON net98 net63 VSS LPNFET W=0.92U L=0.12U M=1 
X17 CON net104 nmcin VSS LPNFET W=0.92U L=0.12U M=1 
X18 net98 B net67 VSS LPNFET W=0.74U L=0.12U M=1 
X19 net98 nmb nma VSS LPNFET W=0.84U L=0.12U M=1 
X2 VDD CI nmcin VDD LPPFET W=1.22U L=0.12U M=1 
X20 net104 B nma VSS LPNFET W=0.88U L=0.12U M=1 
X21 net104 nmb net67 VSS LPNFET W=0.76U L=0.12U M=1 
X3 nmcin CI VSS VSS LPNFET W=0.92U L=0.12U M=1 
X4 VDD B net63 VDD LPPFET W=1.3U L=0.12U M=1 
X5 net63 B VSS VSS LPNFET W=0.92U L=0.12U M=1 
X6 VDD A nma VDD LPPFET W=1.3U L=0.12U M=1 
X7 nma A VSS VSS LPNFET W=0.92U L=0.12U M=1 
X8 VDD nma net67 VDD LPPFET W=1.02U L=0.12U M=1 
X9 net67 nma VSS VSS LPNFET W=0.74U L=0.12U M=1 
.ENDS ACHCONX2TS 

**** 
*.SUBCKT ACHCONX4TS CON A B CI 
.SUBCKT ACHCONX4TS CON A B CI VSS VDD
X0 VDD B net60 VDD LPPFET W=1.3U L=0.12U M=1 
X1 net60 B VSS VSS LPNFET W=0.92U L=0.12U M=1 
X10 CON net105 net64 VDD LPPFET W=1.3U L=0.12U M=1 
X11 CON net99 net62 VDD LPPFET W=2.36U L=0.12U M=1 
X12 net99 net60 net68 VDD LPPFET W=1.24U L=0.12U M=1 
X13 net99 B net66 VDD LPPFET W=1.3U L=0.12U M=1 
X14 net105 net60 net66 VDD LPPFET W=1.28U L=0.12U M=1 
X15 net105 B net68 VDD LPPFET W=1.28U L=0.12U M=1 
X16 CON net99 net64 VSS LPNFET W=0.92U L=0.12U M=1 
X17 CON net105 net62 VSS LPNFET W=1.84U L=0.12U M=1 
X18 net99 B net68 VSS LPNFET W=0.92U L=0.12U M=1 
X19 net99 net60 net66 VSS LPNFET W=0.88U L=0.12U M=1 
X2 VDD CI net62 VDD LPPFET W=2.36U L=0.12U M=1 
X20 net105 B net66 VSS LPNFET W=0.86U L=0.12U M=1 
X21 net105 net60 net68 VSS LPNFET W=0.92U L=0.12U M=1 
X3 net62 CI VSS VSS LPNFET W=1.84U L=0.12U M=1 
X4 VDD B net64 VDD LPPFET W=1.3U L=0.12U M=1 
X5 net64 B VSS VSS LPNFET W=0.92U L=0.12U M=1 
X6 VDD A net66 VDD LPPFET W=1.3U L=0.12U M=1 
X7 net66 A VSS VSS LPNFET W=0.92U L=0.12U M=1 
X8 VDD net66 net68 VDD LPPFET W=1.24U L=0.12U M=1 
X9 net68 net66 VSS VSS LPNFET W=0.92U L=0.12U M=1 
.ENDS ACHCONX4TS 

**** 
*.SUBCKT ADDFHX1TS CO S A B CI 
.SUBCKT ADDFHX1TS CO S A B CI VSS VDD
X0 net103 net121 nmb VDD LPPFET W=0.5U L=0.12U M=1 
X1 net103 net115 nmcin VDD LPPFET W=0.5U L=0.12U M=1 
X10 net109 net115 nmcin VSS LPNFET W=0.36U L=0.12U M=1 
X11 net109 net121 net122 VSS LPNFET W=0.36U L=0.12U M=1 
X12 net115 B net134 VSS LPNFET W=0.52U L=0.12U M=1 
X13 net115 nmb nma VSS LPNFET W=0.52U L=0.12U M=1 
X14 net121 B nma VSS LPNFET W=0.52U L=0.12U M=1 
X15 net121 nmb net134 VSS LPNFET W=0.52U L=0.12U M=1 
X16 VDD nmcin net122 VDD LPPFET W=0.5U L=0.12U M=1 
X17 net122 nmcin VSS VSS LPNFET W=0.36U L=0.12U M=1 
X18 VDD net103 CO VDD LPPFET W=0.64U L=0.12U M=1 
X19 CO net103 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X2 net109 net121 nmcin VDD LPPFET W=0.5U L=0.12U M=1 
X20 VDD net109 S VDD LPPFET W=0.64U L=0.12U M=1 
X21 S net109 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X22 VDD CI nmcin VDD LPPFET W=0.72U L=0.12U M=1 
X23 nmcin CI VSS VSS LPNFET W=0.52U L=0.12U M=1 
X24 VDD B nmb VDD LPPFET W=1.14U L=0.12U M=1 
X25 nmb B VSS VSS LPNFET W=0.82U L=0.12U M=1 
X26 VDD A net132 VDD LPPFET W=0.32U L=0.12U M=1 
X27 net132 A VSS VSS LPNFET W=0.24U L=0.12U M=1 
X28 VDD net132 net134 VDD LPPFET W=0.76U L=0.12U M=1 
X29 net134 net132 VSS VSS LPNFET W=0.52U L=0.12U M=1 
X3 net109 net115 net122 VDD LPPFET W=0.5U L=0.12U M=1 
X30 VDD A nma VDD LPPFET W=0.8U L=0.12U M=1 
X31 nma A VSS VSS LPNFET W=0.58U L=0.12U M=1 
X4 net115 nmb net134 VDD LPPFET W=0.72U L=0.12U M=1 
X5 net115 B nma VDD LPPFET W=0.72U L=0.12U M=1 
X6 net121 nmb nma VDD LPPFET W=0.72U L=0.12U M=1 
X7 net121 B net134 VDD LPPFET W=0.72U L=0.12U M=1 
X8 net103 net115 nmb VSS LPNFET W=0.36U L=0.12U M=1 
X9 net103 net121 nmcin VSS LPNFET W=0.36U L=0.12U M=1 
.ENDS ADDFHX1TS 

**** 
*.SUBCKT ADDFHX2TS CO S A B CI 
.SUBCKT ADDFHX2TS CO S A B CI VSS VDD
X0 net104 net122 nmb VDD LPPFET W=0.96U L=0.12U M=1 
X1 net104 net92 nmcin VDD LPPFET W=0.94U L=0.12U M=1 
X10 net110 net92 nmcin VSS LPNFET W=0.6U L=0.12U M=1 
X11 net110 net122 net123 VSS LPNFET W=0.6U L=0.12U M=1 
X12 net92 B net135 VSS LPNFET W=1.1U L=0.12U M=1 
X13 net92 nmb nma VSS LPNFET W=1.1U L=0.12U M=1 
X14 net122 B nma VSS LPNFET W=1.1U L=0.12U M=1 
X15 net122 nmb net135 VSS LPNFET W=1.1U L=0.12U M=1 
X16 VDD nmcin net123 VDD LPPFET W=1.02U L=0.12U M=1 
X17 net123 nmcin VSS VSS LPNFET W=0.66U L=0.12U M=1 
X18 VDD net104 CO VDD LPPFET W=1.28U L=0.12U M=1 
X19 CO net104 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X2 net110 net122 nmcin VDD LPPFET W=0.92U L=0.12U M=1 
X20 VDD net110 S VDD LPPFET W=1.28U L=0.12U M=1 
X21 S net110 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X22 VDD CI nmcin VDD LPPFET W=1.3U L=0.12U M=1 
X23 nmcin CI VSS VSS LPNFET W=0.92U L=0.12U M=1 
X24 VDD B nmb VDD LPPFET W=2.12U L=0.12U M=1 
X25 nmb B VSS VSS LPNFET W=1.52U L=0.12U M=1 
X26 VDD A net133 VDD LPPFET W=0.66U L=0.12U M=1 
X27 net133 A VSS VSS LPNFET W=0.48U L=0.12U M=1 
X28 VDD net133 net135 VDD LPPFET W=1.64U L=0.12U M=1 
X29 net135 net133 VSS VSS LPNFET W=1.06U L=0.12U M=1 
X3 net110 net92 net123 VDD LPPFET W=1.02U L=0.12U M=1 
X30 VDD A nma VDD LPPFET W=1.64U L=0.12U M=1 
X31 nma A VSS VSS LPNFET W=1.18U L=0.12U M=1 
X4 net92 nmb net135 VDD LPPFET W=1.64U L=0.12U M=1 
X5 net92 B nma VDD LPPFET W=1.64U L=0.12U M=1 
X6 net122 nmb nma VDD LPPFET W=1.64U L=0.12U M=1 
X7 net122 B net135 VDD LPPFET W=1.64U L=0.12U M=1 
X8 net104 net92 nmb VSS LPNFET W=0.6U L=0.12U M=1 
X9 net104 net122 nmcin VSS LPNFET W=0.6U L=0.12U M=1 
.ENDS ADDFHX2TS 

**** 
*.SUBCKT ADDFHX4TS CO S A B CI 
.SUBCKT ADDFHX4TS CO S A B CI VSS VDD
X0 net103 net121 nmb VDD LPPFET W=1.86U L=0.12U M=1 
X1 net103 net115 nmcin VDD LPPFET W=1.86U L=0.12U M=1 
X10 net109 net115 nmcin VSS LPNFET W=1.48U L=0.12U M=1 
X11 net109 net121 net122 VSS LPNFET W=1.4U L=0.12U M=1 
X12 net115 B net134 VSS LPNFET W=2.22U L=0.12U M=1 
X13 net115 nmb nma VSS LPNFET W=2.22U L=0.12U M=1 
X14 net121 B nma VSS LPNFET W=2.22U L=0.12U M=1 
X15 net121 nmb net134 VSS LPNFET W=2.22U L=0.12U M=1 
X16 VDD nmcin net122 VDD LPPFET W=1.96U L=0.12U M=1 
X17 net122 nmcin VSS VSS LPNFET W=1.34U L=0.12U M=1 
X18 VDD net103 CO VDD LPPFET W=2.56U L=0.12U M=1 
X19 CO net103 VSS VSS LPNFET W=1.82U L=0.12U M=1 
X2 net109 net121 nmcin VDD LPPFET W=1.86U L=0.12U M=1 
X20 VDD net109 S VDD LPPFET W=2.56U L=0.12U M=1 
X21 S net109 VSS VSS LPNFET W=1.82U L=0.12U M=1 
X22 VDD CI nmcin VDD LPPFET W=2.58U L=0.12U M=1 
X23 nmcin CI VSS VSS LPNFET W=1.84U L=0.12U M=1 
X24 VDD B nmb VDD LPPFET W=4.32U L=0.12U M=1 
X25 nmb B VSS VSS LPNFET W=3.24U L=0.12U M=1 
X26 VDD A net132 VDD LPPFET W=1.3U L=0.12U M=1 
X27 net132 A VSS VSS LPNFET W=0.8U L=0.12U M=1 
X28 VDD net132 net134 VDD LPPFET W=3.24U L=0.12U M=1 
X29 net134 net132 VSS VSS LPNFET W=2.26U L=0.12U M=1 
X3 net109 net115 net122 VDD LPPFET W=1.86U L=0.12U M=1 
X30 VDD A nma VDD LPPFET W=3.24U L=0.12U M=1 
X31 nma A VSS VSS LPNFET W=2.34U L=0.12U M=1 
X4 net115 nmb net134 VDD LPPFET W=3.18U L=0.12U M=1 
X5 net115 B nma VDD LPPFET W=3.18U L=0.12U M=1 
X6 net121 nmb nma VDD LPPFET W=3.18U L=0.12U M=1 
X7 net121 B net134 VDD LPPFET W=3.18U L=0.12U M=1 
X8 net103 net115 nmb VSS LPNFET W=1.48U L=0.12U M=1 
X9 net103 net121 nmcin VSS LPNFET W=1.52U L=0.12U M=1 
.ENDS ADDFHX4TS 

**** 
*.SUBCKT ADDFHXLTS CO S A B CI 
.SUBCKT ADDFHXLTS CO S A B CI VSS VDD
X0 net103 net121 nmb VDD LPPFET W=0.56U L=0.12U M=1 
X1 net103 net115 nmcin VDD LPPFET W=0.56U L=0.12U M=1 
X10 net109 net115 nmcin VSS LPNFET W=0.32U L=0.12U M=1 
X11 net109 net121 net122 VSS LPNFET W=0.32U L=0.12U M=1 
X12 net115 B net134 VSS LPNFET W=0.32U L=0.12U M=1 
X13 net115 nmb nma VSS LPNFET W=0.32U L=0.12U M=1 
X14 net121 B nma VSS LPNFET W=0.32U L=0.12U M=1 
X15 net121 nmb net134 VSS LPNFET W=0.32U L=0.12U M=1 
X16 VDD nmcin net122 VDD LPPFET W=0.28U L=0.12U M=1 
X17 net122 nmcin VSS VSS LPNFET W=0.2U L=0.12U M=1 
X18 VDD net103 CO VDD LPPFET W=0.42U L=0.12U M=1 
X19 CO net103 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X2 net109 net121 nmcin VDD LPPFET W=0.56U L=0.12U M=1 
X20 VDD net109 S VDD LPPFET W=0.42U L=0.12U M=1 
X21 S net109 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X22 VDD CI nmcin VDD LPPFET W=0.28U L=0.12U M=1 
X23 nmcin CI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X24 VDD B nmb VDD LPPFET W=0.28U L=0.12U M=1 
X25 nmb B VSS VSS LPNFET W=0.2U L=0.12U M=1 
X26 VDD A net132 VDD LPPFET W=0.28U L=0.12U M=1 
X27 net132 A VSS VSS LPNFET W=0.2U L=0.12U M=1 
X28 VDD net132 net134 VDD LPPFET W=0.28U L=0.12U M=1 
X29 net134 net132 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 net109 net115 net122 VDD LPPFET W=0.56U L=0.12U M=1 
X30 VDD A nma VDD LPPFET W=0.28U L=0.12U M=1 
X31 nma A VSS VSS LPNFET W=0.2U L=0.12U M=1 
X4 net115 nmb net134 VDD LPPFET W=0.56U L=0.12U M=1 
X5 net115 B nma VDD LPPFET W=0.56U L=0.12U M=1 
X6 net121 nmb nma VDD LPPFET W=0.56U L=0.12U M=1 
X7 net121 B net134 VDD LPPFET W=0.56U L=0.12U M=1 
X8 net103 net115 nmb VSS LPNFET W=0.32U L=0.12U M=1 
X9 net103 net121 nmcin VSS LPNFET W=0.32U L=0.12U M=1 
.ENDS ADDFHXLTS 

**** 
*.SUBCKT ADDFX1TS CO S A B CI 
.SUBCKT ADDFX1TS CO S A B CI VSS VDD
X0 xo nmb nma VDD LPPFET W=0.5U L=0.12U M=1 
X1 xn net111 nma VDD LPPFET W=0.5U L=0.12U M=1 
X10 xo nma net111 VSS LPNFET W=0.54U L=0.12U M=1 
X11 xn nma nmb VSS LPNFET W=0.54U L=0.12U M=1 
X12 nmcin xo net80 VSS LPNFET W=0.36U L=0.12U M=1 
X13 net80 xn nmb VSS LPNFET W=0.36U L=0.12U M=1 
X14 net110 nmcin xn VSS LPNFET W=0.36U L=0.12U M=1 
X15 net110 CI xo VSS LPNFET W=0.36U L=0.12U M=1 
X16 VDD nmb net111 VDD LPPFET W=0.9U L=0.12U M=1 
X17 net111 nmb VSS VSS LPNFET W=0.64U L=0.12U M=1 
X18 VDD net110 S VDD LPPFET W=0.64U L=0.12U M=1 
X19 S net110 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X2 xn nma net111 VDD LPPFET W=0.76U L=0.12U M=1 
X20 VDD net80 CO VDD LPPFET W=0.64U L=0.12U M=1 
X21 CO net80 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X22 VDD CI nmcin VDD LPPFET W=0.5U L=0.12U M=1 
X23 nmcin CI VSS VSS LPNFET W=0.36U L=0.12U M=1 
X24 VDD B nmb VDD LPPFET W=1.28U L=0.12U M=1 
X25 nmb B VSS VSS LPNFET W=0.92U L=0.12U M=1 
X26 VDD A nma VDD LPPFET W=1.28U L=0.12U M=1 
X27 nma A VSS VSS LPNFET W=0.92U L=0.12U M=1 
X3 xo nma nmb VDD LPPFET W=0.76U L=0.12U M=1 
X4 nmcin xn net80 VDD LPPFET W=0.5U L=0.12U M=1 
X5 net80 xo nmb VDD LPPFET W=0.5U L=0.12U M=1 
X6 net110 CI xn VDD LPPFET W=0.5U L=0.12U M=1 
X7 net110 nmcin xo VDD LPPFET W=0.5U L=0.12U M=1 
X8 xo net111 nma VSS LPNFET W=0.36U L=0.12U M=1 
X9 xn nmb nma VSS LPNFET W=0.36U L=0.12U M=1 
.ENDS ADDFX1TS 

**** 
*.SUBCKT ADDFX2TS CO S A B CI 
.SUBCKT ADDFX2TS CO S A B CI VSS VDD
X0 xo nmb nma VDD LPPFET W=0.5U L=0.12U M=1 
X1 xn net111 nma VDD LPPFET W=0.5U L=0.12U M=1 
X10 xo nma net111 VSS LPNFET W=0.54U L=0.12U M=1 
X11 xn nma nmb VSS LPNFET W=0.54U L=0.12U M=1 
X12 nmcin xo net80 VSS LPNFET W=0.36U L=0.12U M=1 
X13 net80 xn nmb VSS LPNFET W=0.36U L=0.12U M=1 
X14 net110 nmcin xn VSS LPNFET W=0.36U L=0.12U M=1 
X15 net110 CI xo VSS LPNFET W=0.36U L=0.12U M=1 
X16 VDD nmb net111 VDD LPPFET W=0.9U L=0.12U M=1 
X17 net111 nmb VSS VSS LPNFET W=0.64U L=0.12U M=1 
X18 VDD net110 S VDD LPPFET W=1.28U L=0.12U M=1 
X19 S net110 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X2 xn nma net111 VDD LPPFET W=0.76U L=0.12U M=1 
X20 VDD net80 CO VDD LPPFET W=1.28U L=0.12U M=1 
X21 CO net80 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X22 VDD CI nmcin VDD LPPFET W=0.5U L=0.12U M=1 
X23 nmcin CI VSS VSS LPNFET W=0.36U L=0.12U M=1 
X24 VDD B nmb VDD LPPFET W=1.28U L=0.12U M=1 
X25 nmb B VSS VSS LPNFET W=0.92U L=0.12U M=1 
X26 VDD A nma VDD LPPFET W=1.28U L=0.12U M=1 
X27 nma A VSS VSS LPNFET W=0.92U L=0.12U M=1 
X3 xo nma nmb VDD LPPFET W=0.76U L=0.12U M=1 
X4 nmcin xn net80 VDD LPPFET W=0.5U L=0.12U M=1 
X5 net80 xo nmb VDD LPPFET W=0.5U L=0.12U M=1 
X6 net110 CI xn VDD LPPFET W=0.5U L=0.12U M=1 
X7 net110 nmcin xo VDD LPPFET W=0.5U L=0.12U M=1 
X8 xo net111 nma VSS LPNFET W=0.36U L=0.12U M=1 
X9 xn nmb nma VSS LPNFET W=0.36U L=0.12U M=1 
.ENDS ADDFX2TS 

**** 
*.SUBCKT ADDFX4TS CO S A B CI 
.SUBCKT ADDFX4TS CO S A B CI VSS VDD
X0 xo nmb nma VDD LPPFET W=0.5U L=0.12U M=1 
X1 xn net111 nma VDD LPPFET W=0.5U L=0.12U M=1 
X10 xo nma net111 VSS LPNFET W=0.54U L=0.12U M=1 
X11 xn nma nmb VSS LPNFET W=0.54U L=0.12U M=1 
X12 nmcin xo net80 VSS LPNFET W=0.36U L=0.12U M=1 
X13 net80 xn nmb VSS LPNFET W=0.36U L=0.12U M=1 
X14 net110 nmcin xn VSS LPNFET W=0.36U L=0.12U M=1 
X15 net110 CI xo VSS LPNFET W=0.36U L=0.12U M=1 
X16 VDD nmb net111 VDD LPPFET W=0.9U L=0.12U M=1 
X17 net111 nmb VSS VSS LPNFET W=0.64U L=0.12U M=1 
X18 VDD net110 S VDD LPPFET W=2.56U L=0.12U M=1 
X19 S net110 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X2 xn nma net111 VDD LPPFET W=0.68U L=0.12U M=1 
X20 VDD net80 CO VDD LPPFET W=2.56U L=0.12U M=1 
X21 CO net80 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X22 VDD CI nmcin VDD LPPFET W=0.5U L=0.12U M=1 
X23 nmcin CI VSS VSS LPNFET W=0.36U L=0.12U M=1 
X24 VDD B nmb VDD LPPFET W=1.28U L=0.12U M=1 
X25 nmb B VSS VSS LPNFET W=0.9U L=0.12U M=1 
X26 VDD A nma VDD LPPFET W=1.28U L=0.12U M=1 
X27 nma A VSS VSS LPNFET W=0.92U L=0.12U M=1 
X3 xo nma nmb VDD LPPFET W=0.76U L=0.12U M=1 
X4 nmcin xn net80 VDD LPPFET W=0.5U L=0.12U M=1 
X5 net80 xo nmb VDD LPPFET W=0.5U L=0.12U M=1 
X6 net110 CI xn VDD LPPFET W=0.5U L=0.12U M=1 
X7 net110 nmcin xo VDD LPPFET W=0.5U L=0.12U M=1 
X8 xo net111 nma VSS LPNFET W=0.36U L=0.12U M=1 
X9 xn nmb nma VSS LPNFET W=0.36U L=0.12U M=1 
.ENDS ADDFX4TS 

**** 
*.SUBCKT ADDFXLTS CO S A B CI 
.SUBCKT ADDFXLTS CO S A B CI VSS VDD
X0 xo nmb nma VDD LPPFET W=0.56U L=0.12U M=1 
X1 xn net111 nma VDD LPPFET W=0.56U L=0.12U M=1 
X10 xo nma net111 VSS LPNFET W=0.32U L=0.12U M=1 
X11 xn nma nmb VSS LPNFET W=0.32U L=0.12U M=1 
X12 nmcin xo net80 VSS LPNFET W=0.32U L=0.12U M=1 
X13 net80 xn nmb VSS LPNFET W=0.32U L=0.12U M=1 
X14 net110 nmcin xn VSS LPNFET W=0.32U L=0.12U M=1 
X15 net110 CI xo VSS LPNFET W=0.32U L=0.12U M=1 
X16 VDD nmb net111 VDD LPPFET W=0.56U L=0.12U M=1 
X17 net111 nmb VSS VSS LPNFET W=0.32U L=0.12U M=1 
X18 VDD net110 S VDD LPPFET W=0.42U L=0.12U M=1 
X19 S net110 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X2 xn nma net111 VDD LPPFET W=0.56U L=0.12U M=1 
X20 VDD net80 CO VDD LPPFET W=0.42U L=0.12U M=1 
X21 CO net80 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X22 VDD CI nmcin VDD LPPFET W=0.28U L=0.12U M=1 
X23 nmcin CI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X24 VDD B nmb VDD LPPFET W=0.56U L=0.12U M=1 
X25 nmb B VSS VSS LPNFET W=0.32U L=0.12U M=1 
X26 VDD A nma VDD LPPFET W=0.56U L=0.12U M=1 
X27 nma A VSS VSS LPNFET W=0.32U L=0.12U M=1 
X3 xo nma nmb VDD LPPFET W=0.56U L=0.12U M=1 
X4 nmcin xn net80 VDD LPPFET W=0.56U L=0.12U M=1 
X5 net80 xo nmb VDD LPPFET W=0.56U L=0.12U M=1 
X6 net110 CI xn VDD LPPFET W=0.56U L=0.12U M=1 
X7 net110 nmcin xo VDD LPPFET W=0.56U L=0.12U M=1 
X8 xo net111 nma VSS LPNFET W=0.32U L=0.12U M=1 
X9 xn nmb nma VSS LPNFET W=0.32U L=0.12U M=1 
.ENDS ADDFXLTS 

**** 
*.SUBCKT ADDHX1TS CO S A B 
.SUBCKT ADDHX1TS CO S A B VSS VDD
X0 hnet16 A VSS VSS LPNFET W=0.24U L=0.12U M=1 
X1 net27 B hnet16 VSS LPNFET W=0.24U L=0.12U M=1 
X10 VDD B nmb VDD LPPFET W=0.5U L=0.12U M=1 
X11 nmb B VSS VSS LPNFET W=0.36U L=0.12U M=1 
X12 VDD net46 net45 VDD LPPFET W=1.28U L=0.12U M=1 
X13 net45 net46 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X14 VDD A net46 VDD LPPFET W=1.78U L=0.12U M=1 
X15 net46 A VSS VSS LPNFET W=1.28U L=0.12U M=1 
X2 VDD A net27 VDD LPPFET W=0.28U L=0.12U M=1 
X3 VDD B net27 VDD LPPFET W=0.28U L=0.12U M=1 
X4 S B net45 VDD LPPFET W=1.24U L=0.12U M=1 
X5 S nmb net46 VDD LPPFET W=1.24U L=0.12U M=1 
X6 S nmb net45 VSS LPNFET W=0.92U L=0.12U M=1 
X7 S B net46 VSS LPNFET W=0.92U L=0.12U M=1 
X8 VDD net27 CO VDD LPPFET W=0.64U L=0.12U M=1 
X9 CO net27 VSS VSS LPNFET W=0.46U L=0.12U M=1 
.ENDS ADDHX1TS 

**** 
*.SUBCKT ADDHX2TS CO S A B 
.SUBCKT ADDHX2TS CO S A B VSS VDD
X0 hnet16 A VSS VSS LPNFET W=0.48U L=0.12U M=1 
X1 net27 B hnet16 VSS LPNFET W=0.48U L=0.12U M=1 
X10 VDD B nmb VDD LPPFET W=1U L=0.12U M=1 
X11 nmb B VSS VSS LPNFET W=0.74U L=0.12U M=1 
X12 VDD net46 net45 VDD LPPFET W=2.56U L=0.12U M=1 
X13 net45 net46 VSS VSS LPNFET W=1.78U L=0.12U M=1 
X14 VDD A net46 VDD LPPFET W=3.6U L=0.12U M=1 
X15 net46 A VSS VSS LPNFET W=2.58U L=0.12U M=1 
X2 VDD A net27 VDD LPPFET W=0.5U L=0.12U M=1 
X3 VDD B net27 VDD LPPFET W=0.5U L=0.12U M=1 
X4 S B net45 VDD LPPFET W=2.54U L=0.12U M=1 
X5 S nmb net46 VDD LPPFET W=2.54U L=0.12U M=1 
X6 S nmb net45 VSS LPNFET W=1.72U L=0.12U M=1 
X7 S B net46 VSS LPNFET W=1.78U L=0.12U M=1 
X8 VDD net27 CO VDD LPPFET W=1.28U L=0.12U M=1 
X9 CO net27 VSS VSS LPNFET W=0.92U L=0.12U M=1 
.ENDS ADDHX2TS 

**** 
*.SUBCKT ADDHX4TS CO S A B 
.SUBCKT ADDHX4TS CO S A B VSS VDD
X0 hnet16 A VSS VSS LPNFET W=0.92U L=0.12U M=1 
X1 net27 B hnet16 VSS LPNFET W=0.92U L=0.12U M=1 
X10 VDD B nmb VDD LPPFET W=1.96U L=0.12U M=1 
X11 nmb B VSS VSS LPNFET W=1.44U L=0.12U M=1 
X12 VDD net46 net45 VDD LPPFET W=5.12U L=0.12U M=1 
X13 net45 net46 VSS VSS LPNFET W=3.68U L=0.12U M=1 
X14 VDD A net46 VDD LPPFET W=7.18U L=0.12U M=1 
X15 net46 A VSS VSS LPNFET W=4.6U L=0.12U M=1 
X2 VDD A net27 VDD LPPFET W=0.92U L=0.12U M=1 
X3 VDD B net27 VDD LPPFET W=0.92U L=0.12U M=1 
X4 S B net45 VDD LPPFET W=4.96U L=0.12U M=1 
X5 S nmb net46 VDD LPPFET W=4.96U L=0.12U M=1 
X6 S nmb net45 VSS LPNFET W=3.68U L=0.12U M=1 
X7 S B net46 VSS LPNFET W=3.68U L=0.12U M=1 
X8 VDD net27 CO VDD LPPFET W=2.56U L=0.12U M=1 
X9 CO net27 VSS VSS LPNFET W=1.84U L=0.12U M=1 
.ENDS ADDHX4TS 

**** 
*.SUBCKT ADDHXLTS CO S A B 
.SUBCKT ADDHXLTS CO S A B VSS VDD
X0 hnet16 A VSS VSS LPNFET W=0.26U L=0.12U M=1 
X1 net27 B hnet16 VSS LPNFET W=0.26U L=0.12U M=1 
X10 VDD B nmb VDD LPPFET W=0.28U L=0.12U M=1 
X11 nmb B VSS VSS LPNFET W=0.2U L=0.12U M=1 
X12 VDD net46 net45 VDD LPPFET W=0.42U L=0.12U M=1 
X13 net45 net46 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X14 VDD A net46 VDD LPPFET W=0.42U L=0.12U M=1 
X15 net46 A VSS VSS LPNFET W=0.24U L=0.12U M=1 
X2 VDD A net27 VDD LPPFET W=0.28U L=0.12U M=1 
X3 VDD B net27 VDD LPPFET W=0.28U L=0.12U M=1 
X4 S B net45 VDD LPPFET W=0.56U L=0.12U M=1 
X5 S nmb net46 VDD LPPFET W=0.56U L=0.12U M=1 
X6 S nmb net45 VSS LPNFET W=0.32U L=0.12U M=1 
X7 S B net46 VSS LPNFET W=0.32U L=0.12U M=1 
X8 VDD net27 CO VDD LPPFET W=0.42U L=0.12U M=1 
X9 CO net27 VSS VSS LPNFET W=0.24U L=0.12U M=1 
.ENDS ADDHXLTS 

**** 
*.SUBCKT AFCSHCINX2TS CO0 CO1 S A B CI0N CI1N CS 
.SUBCKT AFCSHCINX2TS CO0 CO1 S A B CI0N CI1N CS VSS VDD
X0 net178 CS net233 VDD LPPFET W=0.96U L=0.12U M=1 
X1 net178 net134 net227 VDD LPPFET W=1.02U L=0.12U M=1 
X10 net208 net237 net241 VDD LPPFET W=1.22U L=0.12U M=1 
X11 net208 B net239 VDD LPPFET W=0.98U L=0.12U M=1 
X12 net214 net237 net239 VDD LPPFET W=0.9U L=0.12U M=1 
X13 net214 B net241 VDD LPPFET W=1.22U L=0.12U M=1 
X14 net178 net134 net233 VSS LPNFET W=0.66U L=0.12U M=1 
X15 net178 CS net227 VSS LPNFET W=0.74U L=0.12U M=1 
X16 CO1 net208 net243 VSS LPNFET W=0.6U L=0.12U M=1 
X17 CO1 net214 net229 VSS LPNFET W=0.82U L=0.12U M=1 
X18 net190 net208 net229 VSS LPNFET W=0.58U L=0.12U M=1 
X19 net190 net214 net225 VSS LPNFET W=0.58U L=0.12U M=1 
X2 CO1 net214 net243 VDD LPPFET W=0.98U L=0.12U M=1 
X20 CO0 net208 net219 VSS LPNFET W=0.6U L=0.12U M=1 
X21 CO0 net214 net235 VSS LPNFET W=0.68U L=0.12U M=1 
X22 net202 net208 net235 VSS LPNFET W=0.58U L=0.12U M=1 
X23 net202 net214 net231 VSS LPNFET W=0.58U L=0.12U M=1 
X24 net208 B net241 VSS LPNFET W=0.84U L=0.12U M=1 
X25 net208 net237 net239 VSS LPNFET W=0.66U L=0.12U M=1 
X26 net214 B net239 VSS LPNFET W=0.92U L=0.12U M=1 
X27 net214 net237 net241 VSS LPNFET W=0.58U L=0.12U M=1 
X28 VDD CI1N net215 VDD LPPFET W=0.34U L=0.12U M=1 
X29 net215 CI1N VSS VSS LPNFET W=0.24U L=0.12U M=1 
X3 CO1 net208 net229 VDD LPPFET W=1.3U L=0.12U M=1 
X30 VDD CI0N net217 VDD LPPFET W=0.34U L=0.12U M=1 
X31 net217 CI0N VSS VSS LPNFET W=0.24U L=0.12U M=1 
X32 VDD net237 net219 VDD LPPFET W=1.3U L=0.12U M=1 
X33 net219 net237 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X34 VDD CS net134 VDD LPPFET W=0.42U L=0.12U M=1 
X35 net134 CS VSS VSS LPNFET W=0.3U L=0.12U M=1 
X36 VDD net178 S VDD LPPFET W=1.24U L=0.12U M=1 
X37 S net178 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X38 VDD net215 net225 VDD LPPFET W=0.72U L=0.12U M=1 
X39 net225 net215 VSS VSS LPNFET W=0.58U L=0.12U M=1 
X4 net190 net214 net229 VDD LPPFET W=0.72U L=0.12U M=1 
X40 VDD net190 net227 VDD LPPFET W=1.02U L=0.12U M=1 
X41 net227 net190 VSS VSS LPNFET W=0.74U L=0.12U M=1 
X42 VDD CI1N net229 VDD LPPFET W=1.16U L=0.12U M=1 
X43 net229 CI1N VSS VSS LPNFET W=0.78U L=0.12U M=1 
X44 VDD net217 net231 VDD LPPFET W=0.76U L=0.12U M=1 
X45 net231 net217 VSS VSS LPNFET W=0.58U L=0.12U M=1 
X46 VDD net202 net233 VDD LPPFET W=0.9U L=0.12U M=1 
X47 net233 net202 VSS VSS LPNFET W=0.66U L=0.12U M=1 
X48 VDD CI0N net235 VDD LPPFET W=1.3U L=0.12U M=1 
X49 net235 CI0N VSS VSS LPNFET W=0.92U L=0.12U M=1 
X5 net190 net208 net225 VDD LPPFET W=0.72U L=0.12U M=1 
X50 VDD B net237 VDD LPPFET W=1.3U L=0.12U M=1 
X51 net237 B VSS VSS LPNFET W=0.92U L=0.12U M=1 
X52 VDD A net239 VDD LPPFET W=1.3U L=0.12U M=1 
X53 net239 A VSS VSS LPNFET W=0.92U L=0.12U M=1 
X54 VDD net239 net241 VDD LPPFET W=1.22U L=0.12U M=1 
X55 net241 net239 VSS VSS LPNFET W=0.84U L=0.12U M=1 
X56 VDD net239 net243 VDD LPPFET W=1.3U L=0.12U M=1 
X57 net243 net239 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X6 CO0 net214 net219 VDD LPPFET W=0.98U L=0.12U M=1 
X7 CO0 net208 net235 VDD LPPFET W=1.3U L=0.12U M=1 
X8 net202 net214 net235 VDD LPPFET W=0.8U L=0.12U M=1 
X9 net202 net208 net231 VDD LPPFET W=0.8U L=0.12U M=1 
.ENDS AFCSHCINX2TS 

**** 
*.SUBCKT AFCSHCINX4TS CO0 CO1 S A B CI0N CI1N CS 
.SUBCKT AFCSHCINX4TS CO0 CO1 S A B CI0N CI1N CS VSS VDD
X0 net178 CS net233 VDD LPPFET W=1U L=0.12U M=1 
X1 net178 net134 net227 VDD LPPFET W=1.1U L=0.12U M=1 
X10 net208 net237 net241 VDD LPPFET W=1.28U L=0.12U M=1 
X11 net208 B net239 VDD LPPFET W=0.96U L=0.12U M=1 
X12 net214 net237 net239 VDD LPPFET W=0.92U L=0.12U M=1 
X13 net214 B net241 VDD LPPFET W=1.22U L=0.12U M=1 
X14 net178 net134 net233 VSS LPNFET W=0.6U L=0.12U M=1 
X15 net178 CS net227 VSS LPNFET W=0.58U L=0.12U M=1 
X16 CO1 net208 net243 VSS LPNFET W=1.86U L=0.12U M=1 
X17 CO1 net214 net229 VSS LPNFET W=1.6U L=0.12U M=1 
X18 net190 net208 net229 VSS LPNFET W=0.46U L=0.12U M=1 
X19 net190 net214 net225 VSS LPNFET W=0.46U L=0.12U M=1 
X2 CO1 net214 net243 VDD LPPFET W=2.4U L=0.12U M=1 
X20 CO0 net208 net219 VSS LPNFET W=1.8U L=0.12U M=1 
X21 CO0 net214 net235 VSS LPNFET W=1.72U L=0.12U M=1 
X22 net202 net208 net235 VSS LPNFET W=0.52U L=0.12U M=1 
X23 net202 net214 net231 VSS LPNFET W=0.52U L=0.12U M=1 
X24 net208 B net241 VSS LPNFET W=0.86U L=0.12U M=1 
X25 net208 net237 net239 VSS LPNFET W=0.58U L=0.12U M=1 
X26 net214 B net239 VSS LPNFET W=0.9U L=0.12U M=1 
X27 net214 net237 net241 VSS LPNFET W=0.58U L=0.12U M=1 
X28 VDD CI1N net215 VDD LPPFET W=0.38U L=0.12U M=1 
X29 net215 CI1N VSS VSS LPNFET W=0.26U L=0.12U M=1 
X3 CO1 net208 net229 VDD LPPFET W=1.74U L=0.12U M=1 
X30 VDD CI0N net217 VDD LPPFET W=0.38U L=0.12U M=1 
X31 net217 CI0N VSS VSS LPNFET W=0.28U L=0.12U M=1 
X32 VDD net237 net219 VDD LPPFET W=1.24U L=0.12U M=1 
X33 net219 net237 VSS VSS LPNFET W=0.82U L=0.12U M=1 
X34 VDD CS net134 VDD LPPFET W=0.38U L=0.12U M=1 
X35 net134 CS VSS VSS LPNFET W=0.26U L=0.12U M=1 
X36 VDD net178 S VDD LPPFET W=1.3U L=0.12U M=1 
X37 S net178 VSS VSS LPNFET W=0.86U L=0.12U M=1 
X38 VDD net215 net225 VDD LPPFET W=0.74U L=0.12U M=1 
X39 net225 net215 VSS VSS LPNFET W=0.52U L=0.12U M=1 
X4 net190 net214 net229 VDD LPPFET W=0.74U L=0.12U M=1 
X40 VDD net190 net227 VDD LPPFET W=1.1U L=0.12U M=1 
X41 net227 net190 VSS VSS LPNFET W=0.76U L=0.12U M=1 
X42 VDD CI1N net229 VDD LPPFET W=2.2U L=0.12U M=1 
X43 net229 CI1N VSS VSS LPNFET W=2.06U L=0.12U M=1 
X44 VDD net217 net231 VDD LPPFET W=0.78U L=0.12U M=1 
X45 net231 net217 VSS VSS LPNFET W=0.52U L=0.12U M=1 
X46 VDD net202 net233 VDD LPPFET W=0.98U L=0.12U M=1 
X47 net233 net202 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X48 VDD CI0N net235 VDD LPPFET W=2.92U L=0.12U M=1 
X49 net235 CI0N VSS VSS LPNFET W=1.8U L=0.12U M=1 
X5 net190 net208 net225 VDD LPPFET W=0.74U L=0.12U M=1 
X50 VDD B net237 VDD LPPFET W=1.24U L=0.12U M=1 
X51 net237 B VSS VSS LPNFET W=0.74U L=0.12U M=1 
X52 VDD A net239 VDD LPPFET W=1.28U L=0.12U M=1 
X53 net239 A VSS VSS LPNFET W=0.84U L=0.12U M=1 
X54 VDD net239 net241 VDD LPPFET W=1.28U L=0.12U M=1 
X55 net241 net239 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X56 VDD net239 net243 VDD LPPFET W=1.28U L=0.12U M=1 
X57 net243 net239 VSS VSS LPNFET W=0.84U L=0.12U M=1 
X6 CO0 net214 net219 VDD LPPFET W=2.76U L=0.12U M=1 
X7 CO0 net208 net235 VDD LPPFET W=2.6U L=0.12U M=1 
X8 net202 net214 net235 VDD LPPFET W=0.66U L=0.12U M=1 
X9 net202 net208 net231 VDD LPPFET W=0.78U L=0.12U M=1 
.ENDS AFCSHCINX4TS 

**** 
*.SUBCKT AFCSHCONX2TS CO0N CO1N S A B CI0 CI1 CS 
.SUBCKT AFCSHCONX2TS CO0N CO1N S A B CI0 CI1 CS VSS VDD
X0 net156 CS net207 VDD LPPFET W=1.02U L=0.12U M=1 
X1 net156 net118 net201 VDD LPPFET W=1.02U L=0.12U M=1 
X10 net186 net211 net215 VDD LPPFET W=1.3U L=0.12U M=1 
X11 net186 B net213 VDD LPPFET W=1.3U L=0.12U M=1 
X12 net156 net118 net207 VSS LPNFET W=0.66U L=0.12U M=1 
X13 net156 CS net201 VSS LPNFET W=0.74U L=0.12U M=1 
X14 CO1N net186 net191 VSS LPNFET W=0.86U L=0.12U M=1 
X15 CO1N net193 net187 VSS LPNFET W=0.86U L=0.12U M=1 
X16 net168 net186 net199 VSS LPNFET W=0.58U L=0.12U M=1 
X17 net168 net193 net203 VSS LPNFET W=0.58U L=0.12U M=1 
X18 CO0N net186 net217 VSS LPNFET W=0.92U L=0.12U M=1 
X19 CO0N net193 net189 VSS LPNFET W=0.92U L=0.12U M=1 
X2 CO1N net193 net191 VDD LPPFET W=1.3U L=0.12U M=1 
X20 net180 net186 net205 VSS LPNFET W=0.58U L=0.12U M=1 
X21 net180 net193 net209 VSS LPNFET W=0.58U L=0.12U M=1 
X22 net186 B net215 VSS LPNFET W=0.88U L=0.12U M=1 
X23 net186 net211 net213 VSS LPNFET W=0.92U L=0.12U M=1 
X24 VDD CI1 net187 VDD LPPFET W=1.16U L=0.12U M=1 
X25 net187 CI1 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X26 VDD CI0 net189 VDD LPPFET W=1.3U L=0.12U M=1 
X27 net189 CI0 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X28 VDD B net191 VDD LPPFET W=1.3U L=0.12U M=1 
X29 net191 B VSS VSS LPNFET W=0.92U L=0.12U M=1 
X3 CO1N net186 net187 VDD LPPFET W=1.18U L=0.12U M=1 
X30 VDD net186 net193 VDD LPPFET W=1.3U L=0.12U M=1 
X31 net193 net186 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X32 VDD CS net118 VDD LPPFET W=0.42U L=0.12U M=1 
X33 net118 CS VSS VSS LPNFET W=0.3U L=0.12U M=1 
X34 VDD net156 S VDD LPPFET W=1.28U L=0.12U M=1 
X35 S net156 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X36 VDD net203 net199 VDD LPPFET W=0.8U L=0.12U M=1 
X37 net199 net203 VSS VSS LPNFET W=0.58U L=0.12U M=1 
X38 VDD net168 net201 VDD LPPFET W=1.02U L=0.12U M=1 
X39 net201 net168 VSS VSS LPNFET W=0.74U L=0.12U M=1 
X4 net168 net193 net199 VDD LPPFET W=0.8U L=0.12U M=1 
X40 VDD CI1 net203 VDD LPPFET W=1.16U L=0.12U M=1 
X41 net203 CI1 VSS VSS LPNFET W=0.84U L=0.12U M=1 
X42 VDD net209 net205 VDD LPPFET W=0.8U L=0.12U M=1 
X43 net205 net209 VSS VSS LPNFET W=0.58U L=0.12U M=1 
X44 VDD net180 net207 VDD LPPFET W=0.92U L=0.12U M=1 
X45 net207 net180 VSS VSS LPNFET W=0.66U L=0.12U M=1 
X46 VDD CI0 net209 VDD LPPFET W=1.26U L=0.12U M=1 
X47 net209 CI0 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X48 VDD B net211 VDD LPPFET W=1.3U L=0.12U M=1 
X49 net211 B VSS VSS LPNFET W=0.92U L=0.12U M=1 
X5 net168 net186 net203 VDD LPPFET W=0.8U L=0.12U M=1 
X50 VDD A net213 VDD LPPFET W=1.3U L=0.12U M=1 
X51 net213 A VSS VSS LPNFET W=0.92U L=0.12U M=1 
X52 VDD net213 net215 VDD LPPFET W=1.3U L=0.12U M=1 
X53 net215 net213 VSS VSS LPNFET W=0.88U L=0.12U M=1 
X54 VDD A net217 VDD LPPFET W=1.3U L=0.12U M=1 
X55 net217 A VSS VSS LPNFET W=0.92U L=0.12U M=1 
X6 CO0N net193 net217 VDD LPPFET W=1.2U L=0.12U M=1 
X7 CO0N net186 net189 VDD LPPFET W=1.3U L=0.12U M=1 
X8 net180 net193 net205 VDD LPPFET W=0.8U L=0.12U M=1 
X9 net180 net186 net209 VDD LPPFET W=0.8U L=0.12U M=1 
.ENDS AFCSHCONX2TS 

**** 
*.SUBCKT AFCSHCONX4TS CO0N CO1N S A B CI0 CI1 CS 
.SUBCKT AFCSHCONX4TS CO0N CO1N S A B CI0 CI1 CS VSS VDD
X0 net156 CS net207 VDD LPPFET W=1.02U L=0.12U M=1 
X1 net156 net118 net201 VDD LPPFET W=1.02U L=0.12U M=1 
X10 net186 net211 net215 VDD LPPFET W=1.12U L=0.12U M=1 
X11 net186 B net213 VDD LPPFET W=1.06U L=0.12U M=1 
X12 net156 net118 net207 VSS LPNFET W=0.6U L=0.12U M=1 
X13 net156 CS net201 VSS LPNFET W=0.74U L=0.12U M=1 
X14 CO1N net186 net191 VSS LPNFET W=0.84U L=0.12U M=1 
X15 CO1N net193 net187 VSS LPNFET W=0.92U L=0.12U M=1 
X16 net168 net186 net199 VSS LPNFET W=0.58U L=0.12U M=1 
X17 net168 net193 net203 VSS LPNFET W=0.58U L=0.12U M=1 
X18 CO0N net186 net217 VSS LPNFET W=0.86U L=0.12U M=1 
X19 CO0N net193 net189 VSS LPNFET W=0.9U L=0.12U M=1 
X2 CO1N net193 net191 VDD LPPFET W=1.3U L=0.12U M=1 
X20 net180 net186 net205 VSS LPNFET W=0.5U L=0.12U M=1 
X21 net180 net193 net209 VSS LPNFET W=0.5U L=0.12U M=1 
X22 net186 B net215 VSS LPNFET W=0.72U L=0.12U M=1 
X23 net186 net211 net213 VSS LPNFET W=0.78U L=0.12U M=1 
X24 VDD CI1 net187 VDD LPPFET W=2.2U L=0.12U M=1 
X25 net187 CI1 VSS VSS LPNFET W=1.48U L=0.12U M=1 
X26 VDD CI0 net189 VDD LPPFET W=2.16U L=0.12U M=1 
X27 net189 CI0 VSS VSS LPNFET W=1.82U L=0.12U M=1 
X28 VDD B net191 VDD LPPFET W=1.3U L=0.12U M=1 
X29 net191 B VSS VSS LPNFET W=0.84U L=0.12U M=1 
X3 CO1N net186 net187 VDD LPPFET W=1.3U L=0.12U M=1 
X30 VDD net186 net193 VDD LPPFET W=1.3U L=0.12U M=1 
X31 net193 net186 VSS VSS LPNFET W=0.84U L=0.12U M=1 
X32 VDD CS net118 VDD LPPFET W=0.38U L=0.12U M=1 
X33 net118 CS VSS VSS LPNFET W=0.3U L=0.12U M=1 
X34 VDD net156 S VDD LPPFET W=1.28U L=0.12U M=1 
X35 S net156 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X36 VDD net203 net199 VDD LPPFET W=0.8U L=0.12U M=1 
X37 net199 net203 VSS VSS LPNFET W=0.58U L=0.12U M=1 
X38 VDD net168 net201 VDD LPPFET W=1.02U L=0.12U M=1 
X39 net201 net168 VSS VSS LPNFET W=0.74U L=0.12U M=1 
X4 net168 net193 net199 VDD LPPFET W=0.78U L=0.12U M=1 
X40 VDD CI1 net203 VDD LPPFET W=2.2U L=0.12U M=1 
X41 net203 CI1 VSS VSS LPNFET W=1.48U L=0.12U M=1 
X42 VDD net209 net205 VDD LPPFET W=0.78U L=0.12U M=1 
X43 net205 net209 VSS VSS LPNFET W=0.5U L=0.12U M=1 
X44 VDD net180 net207 VDD LPPFET W=0.98U L=0.12U M=1 
X45 net207 net180 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X46 VDD CI0 net209 VDD LPPFET W=2.16U L=0.12U M=1 
X47 net209 CI0 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X48 VDD B net211 VDD LPPFET W=1.3U L=0.12U M=1 
X49 net211 B VSS VSS LPNFET W=0.84U L=0.12U M=1 
X5 net168 net186 net203 VDD LPPFET W=0.78U L=0.12U M=1 
X50 VDD A net213 VDD LPPFET W=1.3U L=0.12U M=1 
X51 net213 A VSS VSS LPNFET W=0.92U L=0.12U M=1 
X52 VDD net213 net215 VDD LPPFET W=1.12U L=0.12U M=1 
X53 net215 net213 VSS VSS LPNFET W=0.76U L=0.12U M=1 
X54 VDD A net217 VDD LPPFET W=1.3U L=0.12U M=1 
X55 net217 A VSS VSS LPNFET W=0.92U L=0.12U M=1 
X6 CO0N net193 net217 VDD LPPFET W=1.22U L=0.12U M=1 
X7 CO0N net186 net189 VDD LPPFET W=1.3U L=0.12U M=1 
X8 net180 net193 net205 VDD LPPFET W=0.78U L=0.12U M=1 
X9 net180 net186 net209 VDD LPPFET W=0.78U L=0.12U M=1 
.ENDS AFCSHCONX4TS 

**** 
*.SUBCKT AFCSIHCONX2TS CO0N CO1N S A B CS 
.SUBCKT AFCSIHCONX2TS CO0N CO1N S A B CS VSS VDD
X0 CO1N B VSS VSS LPNFET W=0.72U L=0.12U M=1 
X1 CO1N A VSS VSS LPNFET W=0.72U L=0.12U M=1 
X10 VDD nma net61 VDD LPPFET W=0.8U L=0.12U M=1 
X11 net61 nma VSS VSS LPNFET W=0.52U L=0.12U M=1 
X12 VDD net88 S VDD LPPFET W=1.3U L=0.12U M=1 
X13 S net88 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X14 VDD CS nmsel VDD LPPFET W=0.42U L=0.12U M=1 
X15 nmsel CS VSS VSS LPNFET W=0.3U L=0.12U M=1 
X16 VDD B nmb VDD LPPFET W=0.38U L=0.12U M=1 
X17 nmb B VSS VSS LPNFET W=0.28U L=0.12U M=1 
X18 VDD A nma VDD LPPFET W=1.04U L=0.12U M=1 
X19 nma A VSS VSS LPNFET W=0.8U L=0.12U M=1 
X2 VDD B hnet17 VDD LPPFET W=1.3U L=0.12U M=1 
X20 net88 CS net59 VDD LPPFET W=1.02U L=0.12U M=1 
X21 net88 nmsel net94 VDD LPPFET W=0.96U L=0.12U M=1 
X22 net94 nmb nma VDD LPPFET W=1.04U L=0.12U M=1 
X23 net94 B net61 VDD LPPFET W=0.72U L=0.12U M=1 
X24 net88 nmsel net59 VSS LPNFET W=0.74U L=0.12U M=1 
X25 net88 CS net94 VSS LPNFET W=0.74U L=0.12U M=1 
X26 net94 B nma VSS LPNFET W=0.8U L=0.12U M=1 
X27 net94 nmb net61 VSS LPNFET W=0.52U L=0.12U M=1 
X3 hnet17 A CO1N VDD LPPFET W=1.3U L=0.12U M=1 
X4 hnet25 B VSS VSS LPNFET W=0.82U L=0.12U M=1 
X5 CO0N A hnet25 VSS LPNFET W=0.82U L=0.12U M=1 
X6 VDD B CO0N VDD LPPFET W=0.96U L=0.12U M=1 
X7 VDD A CO0N VDD LPPFET W=0.96U L=0.12U M=1 
X8 VDD net94 net59 VDD LPPFET W=1.02U L=0.12U M=1 
X9 net59 net94 VSS VSS LPNFET W=0.74U L=0.12U M=1 
.ENDS AFCSIHCONX2TS 

**** 
*.SUBCKT AFCSIHCONX4TS CO0N CO1N S A B CS 
.SUBCKT AFCSIHCONX4TS CO0N CO1N S A B CS VSS VDD
X0 CO1N B VSS VSS LPNFET W=1.42U L=0.12U M=1 
X1 CO1N A VSS VSS LPNFET W=1.42U L=0.12U M=1 
X10 VDD B CO0N VDD LPPFET W=1.94U L=0.12U M=1 
X11 VDD A CO0N VDD LPPFET W=1.94U L=0.12U M=1 
X12 VDD net94 net59 VDD LPPFET W=1.02U L=0.12U M=1 
X13 net59 net94 VSS VSS LPNFET W=0.74U L=0.12U M=1 
X14 VDD nma net61 VDD LPPFET W=0.8U L=0.12U M=1 
X15 net61 nma VSS VSS LPNFET W=0.52U L=0.12U M=1 
X16 VDD net88 S VDD LPPFET W=1.3U L=0.12U M=1 
X17 S net88 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X18 VDD CS nmsel VDD LPPFET W=0.42U L=0.12U M=1 
X19 nmsel CS VSS VSS LPNFET W=0.3U L=0.12U M=1 
X2 VDD B hnet18 VDD LPPFET W=1.3U L=0.12U M=1 
X20 VDD B nmb VDD LPPFET W=0.38U L=0.12U M=1 
X21 nmb B VSS VSS LPNFET W=0.28U L=0.12U M=1 
X22 VDD A nma VDD LPPFET W=1.04U L=0.12U M=1 
X23 nma A VSS VSS LPNFET W=0.8U L=0.12U M=1 
X24 net88 CS net59 VDD LPPFET W=1.02U L=0.12U M=1 
X25 net88 nmsel net94 VDD LPPFET W=0.96U L=0.12U M=1 
X26 net94 nmb nma VDD LPPFET W=1.04U L=0.12U M=1 
X27 net94 B net61 VDD LPPFET W=0.72U L=0.12U M=1 
X28 net88 nmsel net59 VSS LPNFET W=0.74U L=0.12U M=1 
X29 net88 CS net94 VSS LPNFET W=0.74U L=0.12U M=1 
X3 hnet18 A CO1N VDD LPPFET W=1.3U L=0.12U M=1 
X30 net94 B nma VSS LPNFET W=0.8U L=0.12U M=1 
X31 net94 nmb net61 VSS LPNFET W=0.52U L=0.12U M=1 
X4 VDD B hnet16 VDD LPPFET W=1.3U L=0.12U M=1 
X5 hnet16 A CO1N VDD LPPFET W=1.3U L=0.12U M=1 
X6 hnet27 B VSS VSS LPNFET W=0.82U L=0.12U M=1 
X7 CO0N A hnet27 VSS LPNFET W=0.82U L=0.12U M=1 
X8 hnet23 B VSS VSS LPNFET W=0.82U L=0.12U M=1 
X9 CO0N A hnet23 VSS LPNFET W=0.82U L=0.12U M=1 
.ENDS AFCSIHCONX4TS 

**** 
*.SUBCKT AFHCINX2TS CO S A B CIN 
.SUBCKT AFHCINX2TS CO S A B CIN VSS VDD
X0 VDD CIN net75 VDD LPPFET W=1.3U L=0.12U M=1 
X1 net75 CIN VSS VSS LPNFET W=0.92U L=0.12U M=1 
X10 VDD B net85 VDD LPPFET W=1.12U L=0.12U M=1 
X11 net85 B VSS VSS LPNFET W=0.92U L=0.12U M=1 
X12 VDD A net87 VDD LPPFET W=1.24U L=0.12U M=1 
X13 net87 A VSS VSS LPNFET W=0.92U L=0.12U M=1 
X14 VDD net87 net89 VDD LPPFET W=1.24U L=0.12U M=1 
X15 net89 net87 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X16 CO net138 net77 VDD LPPFET W=1.12U L=0.12U M=1 
X17 CO net132 net75 VDD LPPFET W=1.3U L=0.12U M=1 
X18 net126 net138 net79 VDD LPPFET W=1.02U L=0.12U M=1 
X19 net126 net132 net83 VDD LPPFET W=1.3U L=0.12U M=1 
X2 VDD net85 net77 VDD LPPFET W=1.12U L=0.12U M=1 
X20 net132 net85 net89 VDD LPPFET W=1.24U L=0.12U M=1 
X21 net132 B net87 VDD LPPFET W=1.26U L=0.12U M=1 
X22 net138 net85 net87 VDD LPPFET W=1.22U L=0.12U M=1 
X23 net138 B net89 VDD LPPFET W=1.08U L=0.12U M=1 
X24 CO net132 net77 VSS LPNFET W=0.78U L=0.12U M=1 
X25 CO net138 net75 VSS LPNFET W=0.92U L=0.12U M=1 
X26 net126 net132 net79 VSS LPNFET W=0.74U L=0.12U M=1 
X27 net126 net138 net83 VSS LPNFET W=0.92U L=0.12U M=1 
X28 net132 B net89 VSS LPNFET W=0.92U L=0.12U M=1 
X29 net132 net85 net87 VSS LPNFET W=0.92U L=0.12U M=1 
X3 net77 net85 VSS VSS LPNFET W=0.9U L=0.12U M=1 
X30 net138 B net87 VSS LPNFET W=0.92U L=0.12U M=1 
X31 net138 net85 net89 VSS LPNFET W=0.78U L=0.12U M=1 
X4 VDD net83 net79 VDD LPPFET W=1.02U L=0.12U M=1 
X5 net79 net83 VSS VSS LPNFET W=0.74U L=0.12U M=1 
X6 VDD net126 S VDD LPPFET W=1.18U L=0.12U M=1 
X7 S net126 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X8 VDD CIN net83 VDD LPPFET W=1.3U L=0.12U M=1 
X9 net83 CIN VSS VSS LPNFET W=0.92U L=0.12U M=1 
.ENDS AFHCINX2TS 

**** 
*.SUBCKT AFHCINX4TS CO S A B CIN 
.SUBCKT AFHCINX4TS CO S A B CIN VSS VDD
X0 VDD CIN net75 VDD LPPFET W=2.6U L=0.12U M=1 
X1 net75 CIN VSS VSS LPNFET W=1.8U L=0.12U M=1 
X10 VDD B net85 VDD LPPFET W=1.3U L=0.12U M=1 
X11 net85 B VSS VSS LPNFET W=0.92U L=0.12U M=1 
X12 VDD A net87 VDD LPPFET W=1.3U L=0.12U M=1 
X13 net87 A VSS VSS LPNFET W=0.92U L=0.12U M=1 
X14 VDD net87 net89 VDD LPPFET W=1.3U L=0.12U M=1 
X15 net89 net87 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X16 CO net138 net77 VDD LPPFET W=2.6U L=0.12U M=1 
X17 CO net132 net75 VDD LPPFET W=2.58U L=0.12U M=1 
X18 net126 net138 net79 VDD LPPFET W=1.02U L=0.12U M=1 
X19 net126 net132 net83 VDD LPPFET W=2.58U L=0.12U M=1 
X2 VDD net85 net77 VDD LPPFET W=1.3U L=0.12U M=1 
X20 net132 net85 net89 VDD LPPFET W=1.28U L=0.12U M=1 
X21 net132 B net87 VDD LPPFET W=1.3U L=0.12U M=1 
X22 net138 net85 net87 VDD LPPFET W=1.3U L=0.12U M=1 
X23 net138 B net89 VDD LPPFET W=1.3U L=0.12U M=1 
X24 CO net132 net77 VSS LPNFET W=1.8U L=0.12U M=1 
X25 CO net138 net75 VSS LPNFET W=1.7U L=0.12U M=1 
X26 net126 net132 net79 VSS LPNFET W=0.68U L=0.12U M=1 
X27 net126 net138 net83 VSS LPNFET W=1.82U L=0.12U M=1 
X28 net132 B net89 VSS LPNFET W=0.9U L=0.12U M=1 
X29 net132 net85 net87 VSS LPNFET W=0.92U L=0.12U M=1 
X3 net77 net85 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X30 net138 B net87 VSS LPNFET W=0.92U L=0.12U M=1 
X31 net138 net85 net89 VSS LPNFET W=0.8U L=0.12U M=1 
X4 VDD net83 net79 VDD LPPFET W=1.02U L=0.12U M=1 
X5 net79 net83 VSS VSS LPNFET W=0.68U L=0.12U M=1 
X6 VDD net126 S VDD LPPFET W=1.22U L=0.12U M=1 
X7 S net126 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X8 VDD CIN net83 VDD LPPFET W=2.6U L=0.12U M=1 
X9 net83 CIN VSS VSS LPNFET W=1.8U L=0.12U M=1 
.ENDS AFHCINX4TS 

**** 
*.SUBCKT AFHCONX2TS CON S A B CI 
.SUBCKT AFHCONX2TS CON S A B CI VSS VDD
X0 VDD CI net78 VDD LPPFET W=1.3U L=0.12U M=1 
X1 net78 CI VSS VSS LPNFET W=0.92U L=0.12U M=1 
X10 VDD B net88 VDD LPPFET W=1.3U L=0.12U M=1 
X11 net88 B VSS VSS LPNFET W=0.84U L=0.12U M=1 
X12 VDD A net90 VDD LPPFET W=1.3U L=0.12U M=1 
X13 net90 A VSS VSS LPNFET W=0.92U L=0.12U M=1 
X14 VDD net90 net92 VDD LPPFET W=1.3U L=0.12U M=1 
X15 net92 net90 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X16 CON net141 net88 VDD LPPFET W=1.02U L=0.12U M=1 
X17 CON net135 net78 VDD LPPFET W=1.26U L=0.12U M=1 
X18 net129 net141 net86 VDD LPPFET W=1.02U L=0.12U M=1 
X19 net129 net135 net82 VDD LPPFET W=1.02U L=0.12U M=1 
X2 VDD B net80 VDD LPPFET W=1.3U L=0.12U M=1 
X20 net135 net80 net92 VDD LPPFET W=1.3U L=0.12U M=1 
X21 net135 B net90 VDD LPPFET W=1.3U L=0.12U M=1 
X22 net141 net80 net90 VDD LPPFET W=1.1U L=0.12U M=1 
X23 net141 B net92 VDD LPPFET W=1.24U L=0.12U M=1 
X24 CON net135 net88 VSS LPNFET W=0.74U L=0.12U M=1 
X25 CON net141 net78 VSS LPNFET W=0.84U L=0.12U M=1 
X26 net129 net135 net86 VSS LPNFET W=0.74U L=0.12U M=1 
X27 net129 net141 net82 VSS LPNFET W=0.74U L=0.12U M=1 
X28 net135 B net92 VSS LPNFET W=0.92U L=0.12U M=1 
X29 net135 net80 net90 VSS LPNFET W=0.86U L=0.12U M=1 
X3 net80 B VSS VSS LPNFET W=0.84U L=0.12U M=1 
X30 net141 B net90 VSS LPNFET W=0.78U L=0.12U M=1 
X31 net141 net80 net92 VSS LPNFET W=0.92U L=0.12U M=1 
X4 VDD net86 net82 VDD LPPFET W=1.02U L=0.12U M=1 
X5 net82 net86 VSS VSS LPNFET W=0.72U L=0.12U M=1 
X6 VDD net129 S VDD LPPFET W=1.3U L=0.12U M=1 
X7 S net129 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X8 VDD CI net86 VDD LPPFET W=1.3U L=0.12U M=1 
X9 net86 CI VSS VSS LPNFET W=0.92U L=0.12U M=1 
.ENDS AFHCONX2TS 

**** 
*.SUBCKT AFHCONX4TS CON S A B CI 
.SUBCKT AFHCONX4TS CON S A B CI VSS VDD
X0 VDD CI net78 VDD LPPFET W=2.6U L=0.12U M=1 
X1 net78 CI VSS VSS LPNFET W=1.84U L=0.12U M=1 
X10 VDD B net88 VDD LPPFET W=1.3U L=0.12U M=1 
X11 net88 B VSS VSS LPNFET W=0.84U L=0.12U M=1 
X12 VDD A net90 VDD LPPFET W=1.3U L=0.12U M=1 
X13 net90 A VSS VSS LPNFET W=0.92U L=0.12U M=1 
X14 VDD net90 net92 VDD LPPFET W=1.3U L=0.12U M=1 
X15 net92 net90 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X16 CON net141 net88 VDD LPPFET W=1.02U L=0.12U M=1 
X17 CON net135 net78 VDD LPPFET W=2.52U L=0.12U M=1 
X18 net129 net141 net86 VDD LPPFET W=1.02U L=0.12U M=1 
X19 net129 net135 net82 VDD LPPFET W=1.02U L=0.12U M=1 
X2 VDD B net80 VDD LPPFET W=1.3U L=0.12U M=1 
X20 net135 net80 net92 VDD LPPFET W=1.3U L=0.12U M=1 
X21 net135 B net90 VDD LPPFET W=1.3U L=0.12U M=1 
X22 net141 net80 net90 VDD LPPFET W=1.1U L=0.12U M=1 
X23 net141 B net92 VDD LPPFET W=1.24U L=0.12U M=1 
X24 CON net135 net88 VSS LPNFET W=0.74U L=0.12U M=1 
X25 CON net141 net78 VSS LPNFET W=1.76U L=0.12U M=1 
X26 net129 net135 net86 VSS LPNFET W=0.74U L=0.12U M=1 
X27 net129 net141 net82 VSS LPNFET W=0.74U L=0.12U M=1 
X28 net135 B net92 VSS LPNFET W=0.92U L=0.12U M=1 
X29 net135 net80 net90 VSS LPNFET W=0.86U L=0.12U M=1 
X3 net80 B VSS VSS LPNFET W=0.84U L=0.12U M=1 
X30 net141 B net90 VSS LPNFET W=0.78U L=0.12U M=1 
X31 net141 net80 net92 VSS LPNFET W=0.92U L=0.12U M=1 
X4 VDD net86 net82 VDD LPPFET W=1.02U L=0.12U M=1 
X5 net82 net86 VSS VSS LPNFET W=0.72U L=0.12U M=1 
X6 VDD net129 S VDD LPPFET W=1.3U L=0.12U M=1 
X7 S net129 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X8 VDD CI net86 VDD LPPFET W=2.6U L=0.12U M=1 
X9 net86 CI VSS VSS LPNFET W=1.84U L=0.12U M=1 
.ENDS AFHCONX4TS 

**** 
*.SUBCKT AHCSHCINX2TS CO S A CIN CS 
.SUBCKT AHCSHCINX2TS CO S A CIN CS VSS VDD
X0 CO nma VSS VSS LPNFET W=0.72U L=0.12U M=1 
X1 CO CIN VSS VSS LPNFET W=0.72U L=0.12U M=1 
X10 net69 CS net63 VSS LPNFET W=0.68U L=0.12U M=1 
X11 net63 nmcinn net79 VSS LPNFET W=0.6U L=0.12U M=1 
X12 VDD net69 S VDD LPPFET W=1.3U L=0.12U M=1 
X13 S net69 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X14 VDD CS nmsel VDD LPPFET W=0.42U L=0.12U M=1 
X15 nmsel CS VSS VSS LPNFET W=0.3U L=0.12U M=1 
X16 VDD CIN nmcinn VDD LPPFET W=0.48U L=0.12U M=1 
X17 nmcinn CIN VSS VSS LPNFET W=0.34U L=0.12U M=1 
X18 VDD nma net79 VDD LPPFET W=0.98U L=0.12U M=1 
X19 net79 nma VSS VSS LPNFET W=0.6U L=0.12U M=1 
X2 VDD nma hnet15 VDD LPPFET W=1.3U L=0.12U M=1 
X20 VDD A nma VDD LPPFET W=1.3U L=0.12U M=1 
X21 nma A VSS VSS LPNFET W=0.92U L=0.12U M=1 
X3 hnet15 CIN CO VDD LPPFET W=1.3U L=0.12U M=1 
X4 net63 nmcinn nma VDD LPPFET W=1.28U L=0.12U M=1 
X5 net69 CS nma VDD LPPFET W=0.92U L=0.12U M=1 
X6 net69 nmsel net63 VDD LPPFET W=0.98U L=0.12U M=1 
X7 net63 CIN net79 VDD LPPFET W=1.04U L=0.12U M=1 
X8 net63 CIN nma VSS LPNFET W=0.92U L=0.12U M=1 
X9 net69 nmsel nma VSS LPNFET W=0.68U L=0.12U M=1 
.ENDS AHCSHCINX2TS 

**** 
*.SUBCKT AHCSHCINX4TS CO S A CIN CS 
.SUBCKT AHCSHCINX4TS CO S A CIN CS VSS VDD
X0 CO nma VSS VSS LPNFET W=1.42U L=0.12U M=1 
X1 CO CIN VSS VSS LPNFET W=1.42U L=0.12U M=1 
X10 net63 CIN nma VSS LPNFET W=0.92U L=0.12U M=1 
X11 net69 nmsel nma VSS LPNFET W=0.68U L=0.12U M=1 
X12 net69 CS net63 VSS LPNFET W=0.68U L=0.12U M=1 
X13 net63 nmcinn net79 VSS LPNFET W=0.6U L=0.12U M=1 
X14 VDD net69 S VDD LPPFET W=1.3U L=0.12U M=1 
X15 S net69 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X16 VDD CS nmsel VDD LPPFET W=0.42U L=0.12U M=1 
X17 nmsel CS VSS VSS LPNFET W=0.3U L=0.12U M=1 
X18 VDD CIN nmcinn VDD LPPFET W=0.48U L=0.12U M=1 
X19 nmcinn CIN VSS VSS LPNFET W=0.32U L=0.12U M=1 
X2 VDD nma hnet16 VDD LPPFET W=1.3U L=0.12U M=1 
X20 VDD nma net79 VDD LPPFET W=0.98U L=0.12U M=1 
X21 net79 nma VSS VSS LPNFET W=0.6U L=0.12U M=1 
X22 VDD A nma VDD LPPFET W=1.3U L=0.12U M=1 
X23 nma A VSS VSS LPNFET W=0.92U L=0.12U M=1 
X3 hnet16 CIN CO VDD LPPFET W=1.3U L=0.12U M=1 
X4 VDD nma hnet14 VDD LPPFET W=1.3U L=0.12U M=1 
X5 hnet14 CIN CO VDD LPPFET W=1.3U L=0.12U M=1 
X6 net63 nmcinn nma VDD LPPFET W=1.28U L=0.12U M=1 
X7 net69 CS nma VDD LPPFET W=0.92U L=0.12U M=1 
X8 net69 nmsel net63 VDD LPPFET W=0.98U L=0.12U M=1 
X9 net63 CIN net79 VDD LPPFET W=1.04U L=0.12U M=1 
.ENDS AHCSHCINX4TS 

**** 
*.SUBCKT AHCSHCONX2TS CON S A CI CS 
.SUBCKT AHCSHCONX2TS CON S A CI CS VSS VDD
X0 hnet19 A VSS VSS LPNFET W=0.88U L=0.12U M=1 
X1 CON CI hnet19 VSS LPNFET W=0.88U L=0.12U M=1 
X10 net68 CS net62 VSS LPNFET W=0.74U L=0.12U M=1 
X11 net62 CI net78 VSS LPNFET W=0.74U L=0.12U M=1 
X12 VDD net68 S VDD LPPFET W=1.3U L=0.12U M=1 
X13 S net68 VSS VSS LPNFET W=0.88U L=0.12U M=1 
X14 VDD CS nmsel VDD LPPFET W=0.42U L=0.12U M=1 
X15 nmsel CS VSS VSS LPNFET W=0.3U L=0.12U M=1 
X16 VDD CI nmcin VDD LPPFET W=0.44U L=0.12U M=1 
X17 nmcin CI VSS VSS LPNFET W=0.32U L=0.12U M=1 
X18 VDD nma net78 VDD LPPFET W=0.96U L=0.12U M=1 
X19 net78 nma VSS VSS LPNFET W=0.6U L=0.12U M=1 
X2 VDD A CON VDD LPPFET W=0.96U L=0.12U M=1 
X20 VDD A nma VDD LPPFET W=1.24U L=0.12U M=1 
X21 nma A VSS VSS LPNFET W=0.88U L=0.12U M=1 
X3 VDD CI CON VDD LPPFET W=0.96U L=0.12U M=1 
X4 net62 CI nma VDD LPPFET W=1.24U L=0.12U M=1 
X5 net68 CS nma VDD LPPFET W=0.96U L=0.12U M=1 
X6 net68 nmsel net62 VDD LPPFET W=0.98U L=0.12U M=1 
X7 net62 nmcin net78 VDD LPPFET W=0.96U L=0.12U M=1 
X8 net62 nmcin nma VSS LPNFET W=0.88U L=0.12U M=1 
X9 net68 nmsel nma VSS LPNFET W=0.74U L=0.12U M=1 
.ENDS AHCSHCONX2TS 

**** 
*.SUBCKT AHCSHCONX4TS CON S A CI CS 
.SUBCKT AHCSHCONX4TS CON S A CI CS VSS VDD
X0 hnet20 A VSS VSS LPNFET W=0.92U L=0.12U M=1 
X1 CON CI hnet20 VSS LPNFET W=0.92U L=0.12U M=1 
X10 net62 nmcin nma VSS LPNFET W=0.92U L=0.12U M=1 
X11 net68 nmsel nma VSS LPNFET W=0.68U L=0.12U M=1 
X12 net68 CS net62 VSS LPNFET W=0.68U L=0.12U M=1 
X13 net62 CI net78 VSS LPNFET W=0.74U L=0.12U M=1 
X14 VDD net68 S VDD LPPFET W=1.3U L=0.12U M=1 
X15 S net68 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X16 VDD CS nmsel VDD LPPFET W=0.42U L=0.12U M=1 
X17 nmsel CS VSS VSS LPNFET W=0.3U L=0.12U M=1 
X18 VDD CI nmcin VDD LPPFET W=0.44U L=0.12U M=1 
X19 nmcin CI VSS VSS LPNFET W=0.32U L=0.12U M=1 
X2 hnet14 A VSS VSS LPNFET W=0.92U L=0.12U M=1 
X20 VDD nma net78 VDD LPPFET W=0.98U L=0.12U M=1 
X21 net78 nma VSS VSS LPNFET W=0.6U L=0.12U M=1 
X22 VDD A nma VDD LPPFET W=1.28U L=0.12U M=1 
X23 nma A VSS VSS LPNFET W=0.92U L=0.12U M=1 
X3 CON CI hnet14 VSS LPNFET W=0.92U L=0.12U M=1 
X4 VDD A CON VDD LPPFET W=1.94U L=0.12U M=1 
X5 VDD CI CON VDD LPPFET W=1.94U L=0.12U M=1 
X6 net62 CI nma VDD LPPFET W=1.28U L=0.12U M=1 
X7 net68 CS nma VDD LPPFET W=0.92U L=0.12U M=1 
X8 net68 nmsel net62 VDD LPPFET W=0.98U L=0.12U M=1 
X9 net62 nmcin net78 VDD LPPFET W=0.98U L=0.12U M=1 
.ENDS AHCSHCONX4TS 

**** 
*.SUBCKT AHHCINX2TS CO S A CIN 
.SUBCKT AHHCINX2TS CO S A CIN VSS VDD
X0 CO CIN VSS VSS LPNFET W=0.92U L=0.12U M=1 
X1 CO nmai VSS VSS LPNFET W=0.92U L=0.12U M=1 
X10 VDD A nmai VDD LPPFET W=0.62U L=0.12U M=1 
X11 nmai A VSS VSS LPNFET W=0.44U L=0.12U M=1 
X12 VDD CIN nmcinn VDD LPPFET W=0.5U L=0.12U M=1 
X13 nmcinn CIN VSS VSS LPNFET W=0.36U L=0.12U M=1 
X14 VDD nma net43 VDD LPPFET W=1.28U L=0.12U M=1 
X15 net43 nma VSS VSS LPNFET W=0.92U L=0.12U M=1 
X16 VDD A nma VDD LPPFET W=1.28U L=0.12U M=1 
X17 nma A VSS VSS LPNFET W=0.92U L=0.12U M=1 
X2 VDD CIN hnet13 VDD LPPFET W=0.84U L=0.12U M=1 
X3 hnet13 nmai CO VDD LPPFET W=0.84U L=0.12U M=1 
X4 VDD CIN hnet11 VDD LPPFET W=0.84U L=0.12U M=1 
X5 hnet11 nmai CO VDD LPPFET W=0.84U L=0.12U M=1 
X6 S nmcinn net43 VDD LPPFET W=1.24U L=0.12U M=1 
X7 S CIN nma VDD LPPFET W=1.2U L=0.12U M=1 
X8 S CIN net43 VSS LPNFET W=0.92U L=0.12U M=1 
X9 S nmcinn nma VSS LPNFET W=0.92U L=0.12U M=1 
.ENDS AHHCINX2TS 

**** 
*.SUBCKT AHHCINX4TS CO S A CIN 
.SUBCKT AHHCINX4TS CO S A CIN VSS VDD
X0 CO CIN VSS VSS LPNFET W=1.84U L=0.12U M=1 
X1 CO nmai VSS VSS LPNFET W=1.84U L=0.12U M=1 
X10 S CIN net43 VSS LPNFET W=0.9U L=0.12U M=1 
X11 S nmcinn nma VSS LPNFET W=0.9U L=0.12U M=1 
X12 VDD A nmai VDD LPPFET W=1.2U L=0.12U M=1 
X13 nmai A VSS VSS LPNFET W=0.86U L=0.12U M=1 
X14 VDD CIN nmcinn VDD LPPFET W=0.5U L=0.12U M=1 
X15 nmcinn CIN VSS VSS LPNFET W=0.36U L=0.12U M=1 
X16 VDD nma net43 VDD LPPFET W=1.28U L=0.12U M=1 
X17 net43 nma VSS VSS LPNFET W=0.92U L=0.12U M=1 
X18 VDD A nma VDD LPPFET W=1.22U L=0.12U M=1 
X19 nma A VSS VSS LPNFET W=0.9U L=0.12U M=1 
X2 VDD CIN hnet13 VDD LPPFET W=1.12U L=0.12U M=1 
X3 hnet13 nmai CO VDD LPPFET W=1.12U L=0.12U M=1 
X4 VDD CIN hnet11 VDD LPPFET W=1.12U L=0.12U M=1 
X5 hnet11 nmai CO VDD LPPFET W=1.12U L=0.12U M=1 
X6 VDD CIN hnet15 VDD LPPFET W=1.12U L=0.12U M=1 
X7 hnet15 nmai CO VDD LPPFET W=1.12U L=0.12U M=1 
X8 S nmcinn net43 VDD LPPFET W=1.28U L=0.12U M=1 
X9 S CIN nma VDD LPPFET W=1.22U L=0.12U M=1 
.ENDS AHHCINX4TS 

**** 
*.SUBCKT AHHCONX2TS CON S A CI 
.SUBCKT AHHCONX2TS CON S A CI VSS VDD
X0 hnet16 A VSS VSS LPNFET W=0.58U L=0.12U M=1 
X1 CON CI hnet16 VSS LPNFET W=0.58U L=0.12U M=1 
X10 VDD CI nmcin VDD LPPFET W=0.5U L=0.12U M=1 
X11 nmcin CI VSS VSS LPNFET W=0.36U L=0.12U M=1 
X12 VDD nma net42 VDD LPPFET W=1.28U L=0.12U M=1 
X13 net42 nma VSS VSS LPNFET W=0.92U L=0.12U M=1 
X14 VDD A nma VDD LPPFET W=1.26U L=0.12U M=1 
X15 nma A VSS VSS LPNFET W=0.86U L=0.12U M=1 
X2 hnet10 A VSS VSS LPNFET W=0.58U L=0.12U M=1 
X3 CON CI hnet10 VSS LPNFET W=0.58U L=0.12U M=1 
X4 VDD A CON VDD LPPFET W=1.26U L=0.12U M=1 
X5 VDD CI CON VDD LPPFET W=1.26U L=0.12U M=1 
X6 S CI net42 VDD LPPFET W=1.28U L=0.12U M=1 
X7 S nmcin nma VDD LPPFET W=1.28U L=0.12U M=1 
X8 S nmcin net42 VSS LPNFET W=0.86U L=0.12U M=1 
X9 S CI nma VSS LPNFET W=0.86U L=0.12U M=1 
.ENDS AHHCONX2TS 

**** 
*.SUBCKT AHHCONX4TS CON S A CI 
.SUBCKT AHHCONX4TS CON S A CI VSS VDD
X0 hnet18 A VSS VSS LPNFET W=0.56U L=0.12U M=1 
X1 CON CI hnet18 VSS LPNFET W=0.56U L=0.12U M=1 
X10 S CI net42 VDD LPPFET W=1.28U L=0.12U M=1 
X11 S nmcin nma VDD LPPFET W=1.28U L=0.12U M=1 
X12 S nmcin net42 VSS LPNFET W=0.86U L=0.12U M=1 
X13 S CI nma VSS LPNFET W=0.86U L=0.12U M=1 
X14 VDD CI nmcin VDD LPPFET W=0.5U L=0.12U M=1 
X15 nmcin CI VSS VSS LPNFET W=0.36U L=0.12U M=1 
X16 VDD nma net42 VDD LPPFET W=1.28U L=0.12U M=1 
X17 net42 nma VSS VSS LPNFET W=0.92U L=0.12U M=1 
X18 VDD A nma VDD LPPFET W=1.28U L=0.12U M=1 
X19 nma A VSS VSS LPNFET W=0.86U L=0.12U M=1 
X2 hnet11 A VSS VSS LPNFET W=0.56U L=0.12U M=1 
X3 CON CI hnet11 VSS LPNFET W=0.56U L=0.12U M=1 
X4 hnet13 A VSS VSS LPNFET W=0.56U L=0.12U M=1 
X5 CON CI hnet13 VSS LPNFET W=0.56U L=0.12U M=1 
X6 hnet17 A VSS VSS LPNFET W=0.56U L=0.12U M=1 
X7 CON CI hnet17 VSS LPNFET W=0.56U L=0.12U M=1 
X8 VDD A CON VDD LPPFET W=2.56U L=0.12U M=1 
X9 VDD CI CON VDD LPPFET W=2.56U L=0.12U M=1 
.ENDS AHHCONX4TS 

**** 
*.SUBCKT AND2X1TS Y A B 
.SUBCKT AND2X1TS Y A B VSS VDD
X0 VDD net11 Y VDD LPPFET W=0.64U L=0.12U M=1 
X1 Y net11 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X2 hnet14 B VSS VSS LPNFET W=0.24U L=0.12U M=1 
X3 net11 A hnet14 VSS LPNFET W=0.24U L=0.12U M=1 
X4 VDD B net11 VDD LPPFET W=0.28U L=0.12U M=1 
X5 VDD A net11 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS AND2X1TS 

**** 
*.SUBCKT AND2X2TS Y A B 
.SUBCKT AND2X2TS Y A B VSS VDD
X0 VDD net11 Y VDD LPPFET W=1.28U L=0.12U M=1 
X1 Y net11 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X2 hnet14 B VSS VSS LPNFET W=0.48U L=0.12U M=1 
X3 net11 A hnet14 VSS LPNFET W=0.48U L=0.12U M=1 
X4 VDD B net11 VDD LPPFET W=0.5U L=0.12U M=1 
X5 VDD A net11 VDD LPPFET W=0.5U L=0.12U M=1 
.ENDS AND2X2TS 

**** 
*.SUBCKT AND2X4TS Y A B 
.SUBCKT AND2X4TS Y A B VSS VDD
X0 VDD net11 Y VDD LPPFET W=2.56U L=0.12U M=1 
X1 Y net11 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X2 hnet14 B VSS VSS LPNFET W=0.92U L=0.12U M=1 
X3 net11 A hnet14 VSS LPNFET W=0.92U L=0.12U M=1 
X4 VDD B net11 VDD LPPFET W=0.96U L=0.12U M=1 
X5 VDD A net11 VDD LPPFET W=0.96U L=0.12U M=1 
.ENDS AND2X4TS 

**** 
*.SUBCKT AND2X6TS Y A B 
.SUBCKT AND2X6TS Y A B VSS VDD
X0 VDD net11 Y VDD LPPFET W=3.84U L=0.12U M=1 
X1 Y net11 VSS VSS LPNFET W=2.76U L=0.12U M=1 
X2 hnet15 B VSS VSS LPNFET W=0.66U L=0.12U M=1 
X3 net11 A hnet15 VSS LPNFET W=0.66U L=0.12U M=1 
X4 hnet11 B VSS VSS LPNFET W=0.66U L=0.12U M=1 
X5 net11 A hnet11 VSS LPNFET W=0.66U L=0.12U M=1 
X6 VDD B net11 VDD LPPFET W=1.52U L=0.12U M=1 
X7 VDD A net11 VDD LPPFET W=1.52U L=0.12U M=1 
.ENDS AND2X6TS 

**** 
*.SUBCKT AND2X8TS Y A B
.SUBCKT AND2X8TS Y A B VSS VDD
X0 VDD net11 Y VDD LPPFET W=5.12U L=0.12U M=1 
X1 Y net11 VSS VSS LPNFET W=3.42U L=0.12U M=1 
X2 hnet15 B VSS VSS LPNFET W=0.92U L=0.12U M=1 
X3 net11 A hnet15 VSS LPNFET W=0.92U L=0.12U M=1 
X4 hnet11 B VSS VSS LPNFET W=0.92U L=0.12U M=1 
X5 net11 A hnet11 VSS LPNFET W=0.92U L=0.12U M=1 
X6 VDD B net11 VDD LPPFET W=1.94U L=0.12U M=1 
X7 VDD A net11 VDD LPPFET W=1.94U L=0.12U M=1 
.ENDS AND2X8TS 

**** 
*.SUBCKT AND2XLTS A B Y 
.SUBCKT AND2XLTS A B Y VSS VDD
X0 VDD net11 Y VDD LPPFET W=0.42U L=0.12U M=1 
X1 Y net11 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X2 hnet14 B VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 net11 A hnet14 VSS LPNFET W=0.2U L=0.12U M=1 
X4 VDD B net11 VDD LPPFET W=0.28U L=0.12U M=1 
X5 VDD A net11 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS AND2XLTS 

**** 
*.SUBCKT AND3X1TS Y A B C 
.SUBCKT AND3X1TS Y A B C VSS VDD
X0 VDD net14 Y VDD LPPFET W=0.64U L=0.12U M=1 
X1 Y net14 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X2 hnet17 C VSS VSS LPNFET W=0.3U L=0.12U M=1 
X3 hnet12 B hnet17 VSS LPNFET W=0.3U L=0.12U M=1 
X4 net14 A hnet12 VSS LPNFET W=0.3U L=0.12U M=1 
X5 VDD C net14 VDD LPPFET W=0.28U L=0.12U M=1 
X6 VDD B net14 VDD LPPFET W=0.28U L=0.12U M=1 
X7 VDD A net14 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS AND3X1TS 

**** 
*.SUBCKT AND3X2TS Y A B C 
.SUBCKT AND3X2TS Y A B C VSS VDD
X0 VDD net14 Y VDD LPPFET W=1.28U L=0.12U M=1 
X1 Y net14 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X2 hnet17 C VSS VSS LPNFET W=0.58U L=0.12U M=1 
X3 hnet12 B hnet17 VSS LPNFET W=0.58U L=0.12U M=1 
X4 net14 A hnet12 VSS LPNFET W=0.58U L=0.12U M=1 
X5 VDD C net14 VDD LPPFET W=0.5U L=0.12U M=1 
X6 VDD B net14 VDD LPPFET W=0.5U L=0.12U M=1 
X7 VDD A net14 VDD LPPFET W=0.5U L=0.12U M=1 
.ENDS AND3X2TS 

**** 
*.SUBCKT AND3X4TS Y A B C 
.SUBCKT AND3X4TS Y A B C VSS VDD
X0 hnet15 C VSS VSS LPNFET W=0.92U L=0.12U M=1 
X1 hnet8 B hnet15 VSS LPNFET W=0.92U L=0.12U M=1 
X2 net12 A hnet8 VSS LPNFET W=0.92U L=0.12U M=1 
X3 VDD C net12 VDD LPPFET W=1.02U L=0.12U M=1 
X4 VDD B net12 VDD LPPFET W=1.02U L=0.12U M=1 
X5 VDD A net12 VDD LPPFET W=1.02U L=0.12U M=1 
X6 VDD net12 Y VDD LPPFET W=2.56U L=0.12U M=1 
X7 Y net12 VSS VSS LPNFET W=1.7U L=0.12U M=1 
.ENDS AND3X4TS 

**** 
*.SUBCKT AND3X6TS Y A B C 
.SUBCKT AND3X6TS Y A B C VSS VDD
X0 VDD net14 Y VDD LPPFET W=3.84U L=0.12U M=1 
X1 Y net14 VSS VSS LPNFET W=2.76U L=0.12U M=1 
X10 VDD A net14 VDD LPPFET W=1.44U L=0.12U M=1 
X2 hnet18 C VSS VSS LPNFET W=0.8U L=0.12U M=1 
X3 hnet12 B hnet18 VSS LPNFET W=0.8U L=0.12U M=1 
X4 net14 A hnet12 VSS LPNFET W=0.8U L=0.12U M=1 
X5 hnet19 C VSS VSS LPNFET W=0.8U L=0.12U M=1 
X6 hnet14 B hnet19 VSS LPNFET W=0.8U L=0.12U M=1 
X7 net14 A hnet14 VSS LPNFET W=0.8U L=0.12U M=1 
X8 VDD C net14 VDD LPPFET W=1.44U L=0.12U M=1 
X9 VDD B net14 VDD LPPFET W=1.44U L=0.12U M=1 
.ENDS AND3X6TS 

**** 
*.SUBCKT AND3X8TS Y A B C 
.SUBCKT AND3X8TS Y A B C VSS VDD
X0 hnet16 C VSS VSS LPNFET W=0.92U L=0.12U M=1 
X1 hnet8 B hnet16 VSS LPNFET W=0.92U L=0.12U M=1 
X10 Y net12 VSS VSS LPNFET W=3.68U L=0.12U M=1 
X2 net12 A hnet8 VSS LPNFET W=0.92U L=0.12U M=1 
X3 hnet17 C VSS VSS LPNFET W=0.92U L=0.12U M=1 
X4 hnet11 B hnet17 VSS LPNFET W=0.92U L=0.12U M=1 
X5 net12 A hnet11 VSS LPNFET W=0.92U L=0.12U M=1 
X6 VDD C net12 VDD LPPFET W=2.06U L=0.12U M=1 
X7 VDD B net12 VDD LPPFET W=2.06U L=0.12U M=1 
X8 VDD A net12 VDD LPPFET W=2.06U L=0.12U M=1 
X9 VDD net12 Y VDD LPPFET W=4.64U L=0.12U M=1 
.ENDS AND3X8TS 

**** 
*.SUBCKT AND3XLTS Y A B C 
.SUBCKT AND3XLTS Y A B C VSS VDD
X0 VDD net14 Y VDD LPPFET W=0.42U L=0.12U M=1 
X1 Y net14 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X2 hnet17 C VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 hnet12 B hnet17 VSS LPNFET W=0.2U L=0.12U M=1 
X4 net14 A hnet12 VSS LPNFET W=0.2U L=0.12U M=1 
X5 VDD C net14 VDD LPPFET W=0.28U L=0.12U M=1 
X6 VDD B net14 VDD LPPFET W=0.28U L=0.12U M=1 
X7 VDD A net14 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS AND3XLTS 

**** 
*.SUBCKT AND4X1TS Y A B C D 
.SUBCKT AND4X1TS Y A B C D VSS VDD
X0 VDD net17 Y VDD LPPFET W=0.64U L=0.12U M=1 
X1 Y net17 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X2 hnet14 D VSS VSS LPNFET W=0.32U L=0.12U M=1 
X3 hnet13 C hnet14 VSS LPNFET W=0.32U L=0.12U M=1 
X4 hnet15 B hnet13 VSS LPNFET W=0.32U L=0.12U M=1 
X5 net17 A hnet15 VSS LPNFET W=0.32U L=0.12U M=1 
X6 VDD D net17 VDD LPPFET W=0.28U L=0.12U M=1 
X7 VDD C net17 VDD LPPFET W=0.28U L=0.12U M=1 
X8 VDD B net17 VDD LPPFET W=0.28U L=0.12U M=1 
X9 VDD A net17 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS AND4X1TS 

**** 
*.SUBCKT AND4X2TS Y A B C D 
.SUBCKT AND4X2TS Y A B C D VSS VDD
X0 VDD net17 Y VDD LPPFET W=1.28U L=0.12U M=1 
X1 Y net17 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X2 hnet14 D VSS VSS LPNFET W=0.62U L=0.12U M=1 
X3 hnet13 C hnet14 VSS LPNFET W=0.62U L=0.12U M=1 
X4 hnet15 B hnet13 VSS LPNFET W=0.62U L=0.12U M=1 
X5 net17 A hnet15 VSS LPNFET W=0.62U L=0.12U M=1 
X6 VDD D net17 VDD LPPFET W=0.5U L=0.12U M=1 
X7 VDD C net17 VDD LPPFET W=0.5U L=0.12U M=1 
X8 VDD B net17 VDD LPPFET W=0.5U L=0.12U M=1 
X9 VDD A net17 VDD LPPFET W=0.5U L=0.12U M=1 
.ENDS AND4X2TS 

**** 
*.SUBCKT AND4X4TS Y A B C D 
.SUBCKT AND4X4TS Y A B C D VSS VDD
X0 VDD net17 Y VDD LPPFET W=2.56U L=0.12U M=1 
X1 Y net17 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X10 VDD D net17 VDD LPPFET W=1.04U L=0.12U M=1 
X11 VDD C net17 VDD LPPFET W=1.04U L=0.12U M=1 
X12 VDD B net17 VDD LPPFET W=1.04U L=0.12U M=1 
X13 VDD A net17 VDD LPPFET W=1.04U L=0.12U M=1 
X2 hnet13 D VSS VSS LPNFET W=0.6U L=0.12U M=1 
X3 hnet14 C hnet13 VSS LPNFET W=0.6U L=0.12U M=1 
X4 hnet15 B hnet14 VSS LPNFET W=0.6U L=0.12U M=1 
X5 net17 A hnet15 VSS LPNFET W=0.6U L=0.12U M=1 
X6 hnet18 D VSS VSS LPNFET W=0.6U L=0.12U M=1 
X7 hnet22 C hnet18 VSS LPNFET W=0.6U L=0.12U M=1 
X8 hnet17 B hnet22 VSS LPNFET W=0.6U L=0.12U M=1 
X9 net17 A hnet17 VSS LPNFET W=0.6U L=0.12U M=1 
.ENDS AND4X4TS 

**** 
*.SUBCKT AND4X6TS Y A B C D 
.SUBCKT AND4X6TS Y A B C D VSS VDD
X0 VDD net17 Y VDD LPPFET W=3.84U L=0.12U M=1 
X1 Y net17 VSS VSS LPNFET W=2.5U L=0.12U M=1 
X10 VDD D net17 VDD LPPFET W=1.5U L=0.12U M=1 
X11 VDD C net17 VDD LPPFET W=1.5U L=0.12U M=1 
X12 VDD B net17 VDD LPPFET W=1.5U L=0.12U M=1 
X13 VDD A net17 VDD LPPFET W=1.5U L=0.12U M=1 
X2 hnet13 D VSS VSS LPNFET W=0.92U L=0.12U M=1 
X3 hnet14 C hnet13 VSS LPNFET W=0.92U L=0.12U M=1 
X4 hnet15 B hnet14 VSS LPNFET W=0.92U L=0.12U M=1 
X5 net17 A hnet15 VSS LPNFET W=0.92U L=0.12U M=1 
X6 hnet18 D VSS VSS LPNFET W=0.92U L=0.12U M=1 
X7 hnet22 C hnet18 VSS LPNFET W=0.92U L=0.12U M=1 
X8 hnet17 B hnet22 VSS LPNFET W=0.92U L=0.12U M=1 
X9 net17 A hnet17 VSS LPNFET W=0.92U L=0.12U M=1 
.ENDS AND4X6TS 

**** 
*.SUBCKT AND4X8TS Y A B C D 
.SUBCKT AND4X8TS Y A B C D VSS VDD
X0 VDD net17 Y VDD LPPFET W=5.12U L=0.12U M=1 
X1 Y net17 VSS VSS LPNFET W=3.42U L=0.12U M=1 
X10 hnet17 D VSS VSS LPNFET W=0.8U L=0.12U M=1 
X11 hnet15 C hnet17 VSS LPNFET W=0.8U L=0.12U M=1 
X12 hnet22 B hnet15 VSS LPNFET W=0.8U L=0.12U M=1 
X13 net17 A hnet22 VSS LPNFET W=0.8U L=0.12U M=1 
X14 VDD D net17 VDD LPPFET W=1.92U L=0.12U M=1 
X15 VDD C net17 VDD LPPFET W=1.92U L=0.12U M=1 
X16 VDD B net17 VDD LPPFET W=1.92U L=0.12U M=1 
X17 VDD A net17 VDD LPPFET W=1.92U L=0.12U M=1 
X2 hnet26 D VSS VSS LPNFET W=0.8U L=0.12U M=1 
X3 hnet13 C hnet26 VSS LPNFET W=0.8U L=0.12U M=1 
X4 hnet14 B hnet13 VSS LPNFET W=0.8U L=0.12U M=1 
X5 net17 A hnet14 VSS LPNFET W=0.8U L=0.12U M=1 
X6 hnet18 D VSS VSS LPNFET W=0.8U L=0.12U M=1 
X7 hnet24 C hnet18 VSS LPNFET W=0.8U L=0.12U M=1 
X8 hnet23 B hnet24 VSS LPNFET W=0.8U L=0.12U M=1 
X9 net17 A hnet23 VSS LPNFET W=0.8U L=0.12U M=1 
.ENDS AND4X8TS 

**** 
*.SUBCKT AND4XLTS Y A B C D 
.SUBCKT AND4XLTS Y A B C D VSS VDD
X0 VDD net17 Y VDD LPPFET W=0.42U L=0.12U M=1 
X1 Y net17 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X2 hnet14 D VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 hnet13 C hnet14 VSS LPNFET W=0.2U L=0.12U M=1 
X4 hnet15 B hnet13 VSS LPNFET W=0.2U L=0.12U M=1 
X5 net17 A hnet15 VSS LPNFET W=0.2U L=0.12U M=1 
X6 VDD D net17 VDD LPPFET W=0.28U L=0.12U M=1 
X7 VDD C net17 VDD LPPFET W=0.28U L=0.12U M=1 
X8 VDD B net17 VDD LPPFET W=0.28U L=0.12U M=1 
X9 VDD A net17 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS AND4XLTS 

**** 
*.SUBCKT ANTENNATS A 
.SUBCKT ANTENNATS A VSS VDD
D0 VSS A tdndsx area=0.4898P perim=2.82U 
.ENDS ANTENNATS 

**** 
*.SUBCKT AO21X1TS Y A0 A1 B0 
.SUBCKT AO21X1TS Y A0 A1 B0 VSS VDD
X0 VDD nmin Y VDD LPPFET W=0.64U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=0.46U L=0.12U M=1 
X2 hnet16 A1 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X3 nmin A0 hnet16 VSS LPNFET W=0.24U L=0.12U M=1 
X4 nmin B0 net31 VDD LPPFET W=0.34U L=0.12U M=1 
X5 net31 A1 VDD VDD LPPFET W=0.34U L=0.12U M=1 
X6 net31 A0 VDD VDD LPPFET W=0.34U L=0.12U M=1 
X7 nmin B0 VSS VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS AO21X1TS 

**** 
*.SUBCKT AO21X2TS Y A0 A1 B0 
.SUBCKT AO21X2TS Y A0 A1 B0 VSS VDD
X0 VDD nmin Y VDD LPPFET W=1.28U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=0.86U L=0.12U M=1 
X2 hnet16 A1 VSS VSS LPNFET W=0.48U L=0.12U M=1 
X3 nmin A0 hnet16 VSS LPNFET W=0.48U L=0.12U M=1 
X4 nmin B0 net31 VDD LPPFET W=0.66U L=0.12U M=1 
X5 net31 A1 VDD VDD LPPFET W=0.68U L=0.12U M=1 
X6 net31 A0 VDD VDD LPPFET W=0.66U L=0.12U M=1 
X7 nmin B0 VSS VSS LPNFET W=0.36U L=0.12U M=1 
.ENDS AO21X2TS 

**** 
*.SUBCKT AO21X4TS Y A0 A1 B0 
.SUBCKT AO21X4TS Y A0 A1 B0 VSS VDD
X0 VDD nmin Y VDD LPPFET W=2.46U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=1.84U L=0.12U M=1 
X2 hnet16 A1 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X3 nmin A0 hnet16 VSS LPNFET W=0.92U L=0.12U M=1 
X4 nmin B0 net31 VDD LPPFET W=1.3U L=0.12U M=1 
X5 net31 A1 VDD VDD LPPFET W=1.3U L=0.12U M=1 
X6 net31 A0 VDD VDD LPPFET W=1.3U L=0.12U M=1 
X7 nmin B0 VSS VSS LPNFET W=0.72U L=0.12U M=1 
.ENDS AO21X4TS 

**** 
*.SUBCKT AO21XLTS Y A0 A1 B0 
.SUBCKT AO21XLTS Y A0 A1 B0 VSS VDD
X0 VDD nmin Y VDD LPPFET W=0.42U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=0.24U L=0.12U M=1 
X2 hnet16 A1 VSS VSS LPNFET W=0.26U L=0.12U M=1 
X3 nmin A0 hnet16 VSS LPNFET W=0.26U L=0.12U M=1 
X4 nmin B0 net31 VDD LPPFET W=0.3U L=0.12U M=1 
X5 net31 A1 VDD VDD LPPFET W=0.3U L=0.12U M=1 
X6 net31 A0 VDD VDD LPPFET W=0.3U L=0.12U M=1 
X7 nmin B0 VSS VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS AO21XLTS 

**** 
*.SUBCKT AO22X1TS Y A0 A1 B0 B1 
.SUBCKT AO22X1TS Y A0 A1 B0 B1 VSS VDD
X0 VDD nmin Y VDD LPPFET W=0.64U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=0.46U L=0.12U M=1 
X2 hnet17 A1 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X3 nmin A0 hnet17 VSS LPNFET W=0.24U L=0.12U M=1 
X4 hnet21 B1 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X5 nmin B0 hnet21 VSS LPNFET W=0.24U L=0.12U M=1 
X6 net32 B0 VDD VDD LPPFET W=0.34U L=0.12U M=1 
X7 nmin A0 net32 VDD LPPFET W=0.34U L=0.12U M=1 
X8 net32 B1 VDD VDD LPPFET W=0.34U L=0.12U M=1 
X9 nmin A1 net32 VDD LPPFET W=0.34U L=0.12U M=1 
.ENDS AO22X1TS 

**** 
*.SUBCKT AO22X2TS Y A0 A1 B0 B1 
.SUBCKT AO22X2TS Y A0 A1 B0 B1 VSS VDD
X0 VDD nmin Y VDD LPPFET W=1.28U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=0.86U L=0.12U M=1 
X2 hnet17 A1 VSS VSS LPNFET W=0.48U L=0.12U M=1 
X3 nmin A0 hnet17 VSS LPNFET W=0.48U L=0.12U M=1 
X4 hnet21 B1 VSS VSS LPNFET W=0.48U L=0.12U M=1 
X5 nmin B0 hnet21 VSS LPNFET W=0.48U L=0.12U M=1 
X6 net32 B0 VDD VDD LPPFET W=0.68U L=0.12U M=1 
X7 nmin A0 net32 VDD LPPFET W=0.62U L=0.12U M=1 
X8 net32 B1 VDD VDD LPPFET W=0.68U L=0.12U M=1 
X9 nmin A1 net32 VDD LPPFET W=0.62U L=0.12U M=1 
.ENDS AO22X2TS 

**** 
*.SUBCKT AO22X4TS Y A0 A1 B0 B1 
.SUBCKT AO22X4TS Y A0 A1 B0 B1 VSS VDD
X0 VDD nmin Y VDD LPPFET W=2.34U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=1.84U L=0.12U M=1 
X2 hnet17 A1 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X3 nmin A0 hnet17 VSS LPNFET W=0.92U L=0.12U M=1 
X4 hnet21 B1 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X5 nmin B0 hnet21 VSS LPNFET W=0.92U L=0.12U M=1 
X6 net32 B0 VDD VDD LPPFET W=1.3U L=0.12U M=1 
X7 nmin A0 net32 VDD LPPFET W=1.3U L=0.12U M=1 
X8 net32 B1 VDD VDD LPPFET W=1.3U L=0.12U M=1 
X9 nmin A1 net32 VDD LPPFET W=1.3U L=0.12U M=1 
.ENDS AO22X4TS 

**** 
*.SUBCKT AO22XLTS Y A0 A1 B0 B1 
.SUBCKT AO22XLTS Y A0 A1 B0 B1 VSS VDD
X0 VDD nmin Y VDD LPPFET W=0.42U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=0.24U L=0.12U M=1 
X2 hnet17 A1 VSS VSS LPNFET W=0.26U L=0.12U M=1 
X3 nmin A0 hnet17 VSS LPNFET W=0.26U L=0.12U M=1 
X4 hnet21 B1 VSS VSS LPNFET W=0.26U L=0.12U M=1 
X5 nmin B0 hnet21 VSS LPNFET W=0.26U L=0.12U M=1 
X6 net32 B0 VDD VDD LPPFET W=0.3U L=0.12U M=1 
X7 nmin A0 net32 VDD LPPFET W=0.3U L=0.12U M=1 
X8 net32 B1 VDD VDD LPPFET W=0.3U L=0.12U M=1 
X9 nmin A1 net32 VDD LPPFET W=0.3U L=0.12U M=1 
.ENDS AO22XLTS 

**** 
*.SUBCKT AOI211X1TS Y A0 A1 B0 C0 
.SUBCKT AOI211X1TS Y A0 A1 B0 C0 VSS VDD
X0 hnet15 A1 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X1 Y A0 hnet15 VSS LPNFET W=0.6U L=0.12U M=1 
X2 Y B0 net29 VDD LPPFET W=1.02U L=0.12U M=1 
X3 net29 C0 net35 VDD LPPFET W=1.02U L=0.12U M=1 
X4 net35 A1 VDD VDD LPPFET W=1.02U L=0.12U M=1 
X5 net35 A0 VDD VDD LPPFET W=1.02U L=0.12U M=1 
X6 Y C0 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X7 Y B0 VSS VSS LPNFET W=0.46U L=0.12U M=1 
.ENDS AOI211X1TS 

**** 
*.SUBCKT AOI211X2TS Y A0 A1 B0 C0 
.SUBCKT AOI211X2TS Y A0 A1 B0 C0 VSS VDD
X0 hnet17 A1 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X1 Y A0 hnet17 VSS LPNFET W=0.6U L=0.12U M=1 
X10 Y C0 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X11 Y B0 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X2 hnet13 A1 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X3 Y A0 hnet13 VSS LPNFET W=0.6U L=0.12U M=1 
X4 Y B0 net30 VDD LPPFET W=1.04U L=0.12U M=1 
X5 net30 C0 net42 VDD LPPFET W=1.04U L=0.12U M=1 
X6 Y B0 net36 VDD LPPFET W=1.04U L=0.12U M=1 
X7 net36 C0 net42 VDD LPPFET W=1.04U L=0.12U M=1 
X8 net42 A1 VDD VDD LPPFET W=2.06U L=0.12U M=1 
X9 net42 A0 VDD VDD LPPFET W=2.06U L=0.12U M=1 
.ENDS AOI211X2TS 

**** 
*.SUBCKT AOI211X4TS Y A0 A1 B0 C0 
.SUBCKT AOI211X4TS Y A0 A1 B0 C0 VSS VDD
X0 VDD net26 net22 VDD LPPFET W=1.02U L=0.12U M=1 
X1 net22 net26 VSS VSS LPNFET W=0.74U L=0.12U M=1 
X10 net26 C0 VSS VSS LPNFET W=0.3U L=0.12U M=1 
X11 net26 B0 VSS VSS LPNFET W=0.3U L=0.12U M=1 
X2 VDD net22 Y VDD LPPFET W=2.56U L=0.12U M=1 
X3 Y net22 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X4 hnet21 A1 VSS VSS LPNFET W=0.38U L=0.12U M=1 
X5 net26 A0 hnet21 VSS LPNFET W=0.38U L=0.12U M=1 
X6 net26 B0 net34 VDD LPPFET W=0.66U L=0.12U M=1 
X7 net34 C0 net40 VDD LPPFET W=0.66U L=0.12U M=1 
X8 net40 A1 VDD VDD LPPFET W=0.66U L=0.12U M=1 
X9 net40 A0 VDD VDD LPPFET W=0.66U L=0.12U M=1 
.ENDS AOI211X4TS 

**** 
*.SUBCKT AOI211XLTS Y A0 A1 B0 C0 
.SUBCKT AOI211XLTS Y A0 A1 B0 C0 VSS VDD
X0 hnet15 A1 VSS VSS LPNFET W=0.4U L=0.12U M=1 
X1 Y A0 hnet15 VSS LPNFET W=0.4U L=0.12U M=1 
X2 Y B0 net29 VDD LPPFET W=0.54U L=0.12U M=1 
X3 net29 C0 net35 VDD LPPFET W=0.54U L=0.12U M=1 
X4 net35 A1 VDD VDD LPPFET W=0.54U L=0.12U M=1 
X5 net35 A0 VDD VDD LPPFET W=0.54U L=0.12U M=1 
X6 Y C0 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X7 Y B0 VSS VSS LPNFET W=0.24U L=0.12U M=1 
.ENDS AOI211XLTS 

**** 
*.SUBCKT AOI21X1TS Y A0 A1 B0 
.SUBCKT AOI21X1TS Y A0 A1 B0 VSS VDD
X0 hnet13 A1 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X1 Y A0 hnet13 VSS LPNFET W=0.6U L=0.12U M=1 
X2 Y B0 net29 VDD LPPFET W=0.84U L=0.12U M=1 
X3 net29 A1 VDD VDD LPPFET W=0.84U L=0.12U M=1 
X4 net29 A0 VDD VDD LPPFET W=0.84U L=0.12U M=1 
X5 Y B0 VSS VSS LPNFET W=0.46U L=0.12U M=1 
.ENDS AOI21X1TS 

**** 
*.SUBCKT AOI21X2TS Y A0 A1 B0 
.SUBCKT AOI21X2TS Y A0 A1 B0 VSS VDD
X0 hnet14 A1 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X1 Y A0 hnet14 VSS LPNFET W=0.6U L=0.12U M=1 
X2 hnet10 A1 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X3 Y A0 hnet10 VSS LPNFET W=0.6U L=0.12U M=1 
X4 Y B0 net29 VDD LPPFET W=1.68U L=0.12U M=1 
X5 net29 A1 VDD VDD LPPFET W=1.68U L=0.12U M=1 
X6 net29 A0 VDD VDD LPPFET W=1.68U L=0.12U M=1 
X7 Y B0 VSS VSS LPNFET W=0.92U L=0.12U M=1 
.ENDS AOI21X2TS 

**** 
*.SUBCKT AOI21X4TS Y A0 A1 B0 
.SUBCKT AOI21X4TS Y A0 A1 B0 VSS VDD
X0 hnet15 A1 VSS VSS LPNFET W=0.82U L=0.12U M=1 
X1 Y A0 hnet15 VSS LPNFET W=0.82U L=0.12U M=1 
X2 hnet10 A1 VSS VSS LPNFET W=0.82U L=0.12U M=1 
X3 Y A0 hnet10 VSS LPNFET W=0.82U L=0.12U M=1 
X4 hnet14 A1 VSS VSS LPNFET W=0.82U L=0.12U M=1 
X5 Y A0 hnet14 VSS LPNFET W=0.82U L=0.12U M=1 
X6 Y B0 net29 VDD LPPFET W=3.36U L=0.12U M=1 
X7 net29 A1 VDD VDD LPPFET W=3.36U L=0.12U M=1 
X8 net29 A0 VDD VDD LPPFET W=3.36U L=0.12U M=1 
X9 Y B0 VSS VSS LPNFET W=1.84U L=0.12U M=1 
.ENDS AOI21X4TS 

**** 
*.SUBCKT AOI21XLTS Y A0 A1 B0 
.SUBCKT AOI21XLTS Y A0 A1 B0 VSS VDD
X0 hnet13 A1 VSS VSS LPNFET W=0.4U L=0.12U M=1 
X1 Y A0 hnet13 VSS LPNFET W=0.4U L=0.12U M=1 
X2 Y B0 net29 VDD LPPFET W=0.44U L=0.12U M=1 
X3 net29 A1 VDD VDD LPPFET W=0.44U L=0.12U M=1 
X4 net29 A0 VDD VDD LPPFET W=0.44U L=0.12U M=1 
X5 Y B0 VSS VSS LPNFET W=0.24U L=0.12U M=1 
.ENDS AOI21XLTS 

**** 
*.SUBCKT AOI221X1TS Y A0 A1 B0 B1 C0 
.SUBCKT AOI221X1TS Y A0 A1 B0 B1 C0 VSS VDD
X0 hnet16 B1 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X1 Y B0 hnet16 VSS LPNFET W=0.6U L=0.12U M=1 
X2 hnet20 A1 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X3 Y A0 hnet20 VSS LPNFET W=0.6U L=0.12U M=1 
X4 Y C0 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X5 Y C0 net46 VDD LPPFET W=1.02U L=0.12U M=1 
X6 net43 B0 VDD VDD LPPFET W=1.02U L=0.12U M=1 
X7 net46 A0 net43 VDD LPPFET W=1.02U L=0.12U M=1 
X8 net43 B1 VDD VDD LPPFET W=1.02U L=0.12U M=1 
X9 net46 A1 net43 VDD LPPFET W=1.02U L=0.12U M=1 
.ENDS AOI221X1TS 

**** 
*.SUBCKT AOI221X2TS Y A0 A1 B0 B1 C0 
.SUBCKT AOI221X2TS Y A0 A1 B0 B1 C0 VSS VDD
X0 hnet17 B1 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X1 Y B0 hnet17 VSS LPNFET W=0.6U L=0.12U M=1 
X10 net43 B0 VDD VDD LPPFET W=2.06U L=0.12U M=1 
X11 net46 A0 net43 VDD LPPFET W=2.06U L=0.12U M=1 
X12 net43 B1 VDD VDD LPPFET W=2.06U L=0.12U M=1 
X13 net46 A1 net43 VDD LPPFET W=2.06U L=0.12U M=1 
X2 hnet13 B1 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X3 Y B0 hnet13 VSS LPNFET W=0.6U L=0.12U M=1 
X4 hnet22 A1 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X5 Y A0 hnet22 VSS LPNFET W=0.6U L=0.12U M=1 
X6 hnet18 A1 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X7 Y A0 hnet18 VSS LPNFET W=0.6U L=0.12U M=1 
X8 Y C0 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X9 Y C0 net46 VDD LPPFET W=2.06U L=0.12U M=1 
.ENDS AOI221X2TS 

**** 
*.SUBCKT AOI221X4TS Y A0 A1 B0 B1 C0 
.SUBCKT AOI221X4TS Y A0 A1 B0 B1 C0 VSS VDD
X0 VDD nmin net24 VDD LPPFET W=1.02U L=0.12U M=1 
X1 net24 nmin VSS VSS LPNFET W=0.74U L=0.12U M=1 
X10 net48 B0 VDD VDD LPPFET W=0.66U L=0.12U M=1 
X11 net51 A0 net48 VDD LPPFET W=0.66U L=0.12U M=1 
X12 net48 B1 VDD VDD LPPFET W=0.66U L=0.12U M=1 
X13 net51 A1 net48 VDD LPPFET W=0.66U L=0.12U M=1 
X2 VDD net24 Y VDD LPPFET W=2.56U L=0.12U M=1 
X3 Y net24 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X4 hnet22 B1 VSS VSS LPNFET W=0.38U L=0.12U M=1 
X5 nmin B0 hnet22 VSS LPNFET W=0.38U L=0.12U M=1 
X6 hnet26 A1 VSS VSS LPNFET W=0.38U L=0.12U M=1 
X7 nmin A0 hnet26 VSS LPNFET W=0.38U L=0.12U M=1 
X8 nmin C0 VSS VSS LPNFET W=0.3U L=0.12U M=1 
X9 nmin C0 net51 VDD LPPFET W=0.66U L=0.12U M=1 
.ENDS AOI221X4TS 

**** 
*.SUBCKT AOI221XLTS Y A0 A1 B0 B1 C0 
.SUBCKT AOI221XLTS Y A0 A1 B0 B1 C0 VSS VDD
X0 hnet16 B1 VSS VSS LPNFET W=0.4U L=0.12U M=1 
X1 Y B0 hnet16 VSS LPNFET W=0.4U L=0.12U M=1 
X2 hnet20 A1 VSS VSS LPNFET W=0.4U L=0.12U M=1 
X3 Y A0 hnet20 VSS LPNFET W=0.4U L=0.12U M=1 
X4 Y C0 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X5 Y C0 net46 VDD LPPFET W=0.54U L=0.12U M=1 
X6 net43 B0 VDD VDD LPPFET W=0.54U L=0.12U M=1 
X7 net46 A0 net43 VDD LPPFET W=0.54U L=0.12U M=1 
X8 net43 B1 VDD VDD LPPFET W=0.54U L=0.12U M=1 
X9 net46 A1 net43 VDD LPPFET W=0.54U L=0.12U M=1 
.ENDS AOI221XLTS 

**** 
*.SUBCKT AOI222X1TS Y A0 A1 B0 B1 C0 C1 
.SUBCKT AOI222X1TS Y A0 A1 B0 B1 C0 C1 VSS VDD
X0 hnet16 C1 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X1 Y C0 hnet16 VSS LPNFET W=0.6U L=0.12U M=1 
X10 net55 C1 VDD VDD LPPFET W=1.02U L=0.12U M=1 
X11 Y A1 net46 VDD LPPFET W=1.02U L=0.12U M=1 
X2 hnet21 B1 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X3 Y B0 hnet21 VSS LPNFET W=0.6U L=0.12U M=1 
X4 hnet26 A1 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X5 Y A0 hnet26 VSS LPNFET W=0.6U L=0.12U M=1 
X6 net46 B0 net55 VDD LPPFET W=1.02U L=0.12U M=1 
X7 net46 B1 net55 VDD LPPFET W=1.02U L=0.12U M=1 
X8 net55 C0 VDD VDD LPPFET W=1.02U L=0.12U M=1 
X9 Y A0 net46 VDD LPPFET W=1.02U L=0.12U M=1 
.ENDS AOI222X1TS 

**** 
*.SUBCKT AOI222X2TS Y A0 A1 B0 B1 C0 C1 
.SUBCKT AOI222X2TS Y A0 A1 B0 B1 C0 C1 VSS VDD
X0 hnet18 C1 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X1 Y C0 hnet18 VSS LPNFET W=0.6U L=0.12U M=1 
X10 hnet25 A1 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X11 Y A0 hnet25 VSS LPNFET W=0.6U L=0.12U M=1 
X12 net46 B0 net55 VDD LPPFET W=2.06U L=0.12U M=1 
X13 net46 B1 net55 VDD LPPFET W=2.06U L=0.12U M=1 
X14 net55 C0 VDD VDD LPPFET W=2.06U L=0.12U M=1 
X15 Y A0 net46 VDD LPPFET W=2.06U L=0.12U M=1 
X16 net55 C1 VDD VDD LPPFET W=2.06U L=0.12U M=1 
X17 Y A1 net46 VDD LPPFET W=2.06U L=0.12U M=1 
X2 hnet13 C1 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X3 Y C0 hnet13 VSS LPNFET W=0.6U L=0.12U M=1 
X4 hnet24 B1 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X5 Y B0 hnet24 VSS LPNFET W=0.6U L=0.12U M=1 
X6 hnet19 B1 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X7 Y B0 hnet19 VSS LPNFET W=0.6U L=0.12U M=1 
X8 hnet30 A1 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X9 Y A0 hnet30 VSS LPNFET W=0.6U L=0.12U M=1 
.ENDS AOI222X2TS 

**** 
*.SUBCKT AOI222X4TS Y A0 A1 B0 B1 C0 C1 
.SUBCKT AOI222X4TS Y A0 A1 B0 B1 C0 C1 VSS VDD
X0 VDD nmin net33 VDD LPPFET W=1.02U L=0.12U M=1 
X1 net33 nmin VSS VSS LPNFET W=0.74U L=0.12U M=1 
X10 net51 B0 net60 VDD LPPFET W=0.66U L=0.12U M=1 
X11 net51 B1 net60 VDD LPPFET W=0.66U L=0.12U M=1 
X12 net60 C0 VDD VDD LPPFET W=0.66U L=0.12U M=1 
X13 nmin A0 net51 VDD LPPFET W=0.66U L=0.12U M=1 
X14 net60 C1 VDD VDD LPPFET W=0.66U L=0.12U M=1 
X15 nmin A1 net51 VDD LPPFET W=0.66U L=0.12U M=1 
X2 VDD net33 Y VDD LPPFET W=2.56U L=0.12U M=1 
X3 Y net33 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X4 hnet24 C1 VSS VSS LPNFET W=0.38U L=0.12U M=1 
X5 nmin C0 hnet24 VSS LPNFET W=0.38U L=0.12U M=1 
X6 hnet28 B1 VSS VSS LPNFET W=0.38U L=0.12U M=1 
X7 nmin B0 hnet28 VSS LPNFET W=0.38U L=0.12U M=1 
X8 hnet32 A1 VSS VSS LPNFET W=0.38U L=0.12U M=1 
X9 nmin A0 hnet32 VSS LPNFET W=0.38U L=0.12U M=1 
.ENDS AOI222X4TS 

**** 
*.SUBCKT AOI222XLTS Y A0 A1 B0 B1 C0 C1 
.SUBCKT AOI222XLTS Y A0 A1 B0 B1 C0 C1 VSS VDD
X0 hnet16 C1 VSS VSS LPNFET W=0.4U L=0.12U M=1 
X1 Y C0 hnet16 VSS LPNFET W=0.4U L=0.12U M=1 
X10 Y A0 net49 VDD LPPFET W=0.54U L=0.12U M=1 
X11 Y A1 net49 VDD LPPFET W=0.54U L=0.12U M=1 
X2 hnet21 B1 VSS VSS LPNFET W=0.4U L=0.12U M=1 
X3 Y B0 hnet21 VSS LPNFET W=0.4U L=0.12U M=1 
X4 hnet26 A1 VSS VSS LPNFET W=0.4U L=0.12U M=1 
X5 Y A0 hnet26 VSS LPNFET W=0.4U L=0.12U M=1 
X6 net43 C1 VDD VDD LPPFET W=0.54U L=0.12U M=1 
X7 net49 B0 net43 VDD LPPFET W=0.54U L=0.12U M=1 
X8 net49 B1 net43 VDD LPPFET W=0.54U L=0.12U M=1 
X9 net43 C0 VDD VDD LPPFET W=0.54U L=0.12U M=1 
.ENDS AOI222XLTS 

**** 
*.SUBCKT AOI22X1TS Y A0 A1 B0 B1 
.SUBCKT AOI22X1TS Y A0 A1 B0 B1 VSS VDD
X0 hnet13 A1 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X1 Y A0 hnet13 VSS LPNFET W=0.6U L=0.12U M=1 
X2 hnet18 B1 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X3 Y B0 hnet18 VSS LPNFET W=0.6U L=0.12U M=1 
X4 net30 B0 VDD VDD LPPFET W=0.84U L=0.12U M=1 
X5 Y A0 net30 VDD LPPFET W=0.84U L=0.12U M=1 
X6 net30 B1 VDD VDD LPPFET W=0.84U L=0.12U M=1 
X7 Y A1 net30 VDD LPPFET W=0.84U L=0.12U M=1 
.ENDS AOI22X1TS 

**** 
*.SUBCKT AOI22X2TS Y A0 A1 B0 B1 
.SUBCKT AOI22X2TS Y A0 A1 B0 B1 VSS VDD
X0 hnet15 A1 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X1 Y A0 hnet15 VSS LPNFET W=0.6U L=0.12U M=1 
X10 net30 B1 VDD VDD LPPFET W=1.68U L=0.12U M=1 
X11 Y A1 net30 VDD LPPFET W=1.68U L=0.12U M=1 
X2 hnet10 A1 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X3 Y A0 hnet10 VSS LPNFET W=0.6U L=0.12U M=1 
X4 hnet21 B1 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X5 Y B0 hnet21 VSS LPNFET W=0.6U L=0.12U M=1 
X6 hnet16 B1 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X7 Y B0 hnet16 VSS LPNFET W=0.6U L=0.12U M=1 
X8 net30 B0 VDD VDD LPPFET W=1.68U L=0.12U M=1 
X9 Y A0 net30 VDD LPPFET W=1.68U L=0.12U M=1 
.ENDS AOI22X2TS 

**** 
*.SUBCKT AOI22X4TS Y A0 A1 B0 B1 
.SUBCKT AOI22X4TS Y A0 A1 B0 B1 VSS VDD
X0 hnet16 A1 VSS VSS LPNFET W=0.82U L=0.12U M=1 
X1 Y A0 hnet16 VSS LPNFET W=0.82U L=0.12U M=1 
X10 hnet22 B1 VSS VSS LPNFET W=0.82U L=0.12U M=1 
X11 Y B0 hnet22 VSS LPNFET W=0.82U L=0.12U M=1 
X12 net30 B0 VDD VDD LPPFET W=3.36U L=0.12U M=1 
X13 Y A0 net30 VDD LPPFET W=3.36U L=0.12U M=1 
X14 net30 B1 VDD VDD LPPFET W=3.36U L=0.12U M=1 
X15 Y A1 net30 VDD LPPFET W=3.36U L=0.12U M=1 
X2 hnet10 A1 VSS VSS LPNFET W=0.82U L=0.12U M=1 
X3 Y A0 hnet10 VSS LPNFET W=0.82U L=0.12U M=1 
X4 hnet15 A1 VSS VSS LPNFET W=0.82U L=0.12U M=1 
X5 Y A0 hnet15 VSS LPNFET W=0.82U L=0.12U M=1 
X6 hnet23 B1 VSS VSS LPNFET W=0.82U L=0.12U M=1 
X7 Y B0 hnet23 VSS LPNFET W=0.82U L=0.12U M=1 
X8 hnet17 B1 VSS VSS LPNFET W=0.82U L=0.12U M=1 
X9 Y B0 hnet17 VSS LPNFET W=0.82U L=0.12U M=1 
.ENDS AOI22X4TS 

**** 
*.SUBCKT AOI22XLTS Y A0 A1 B0 B1 
.SUBCKT AOI22XLTS Y A0 A1 B0 B1 VSS VDD
X0 hnet13 A1 VSS VSS LPNFET W=0.4U L=0.12U M=1 
X1 Y A0 hnet13 VSS LPNFET W=0.4U L=0.12U M=1 
X2 hnet18 B1 VSS VSS LPNFET W=0.4U L=0.12U M=1 
X3 Y B0 hnet18 VSS LPNFET W=0.4U L=0.12U M=1 
X4 net30 B0 VDD VDD LPPFET W=0.44U L=0.12U M=1 
X5 Y A0 net30 VDD LPPFET W=0.44U L=0.12U M=1 
X6 net30 B1 VDD VDD LPPFET W=0.44U L=0.12U M=1 
X7 Y A1 net30 VDD LPPFET W=0.44U L=0.12U M=1 
.ENDS AOI22XLTS 

**** 
*.SUBCKT AOI2BB1X1TS Y A0N A1N B0 
.SUBCKT AOI2BB1X1TS Y A0N A1N B0 VSS VDD
X0 Y B0 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X1 Y net13 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X2 VDD B0 hnet9 VDD LPPFET W=0.84U L=0.12U M=1 
X3 hnet9 net13 Y VDD LPPFET W=0.84U L=0.12U M=1 
X4 net13 A1N VSS VSS LPNFET W=0.22U L=0.12U M=1 
X5 net13 A0N VSS VSS LPNFET W=0.22U L=0.12U M=1 
X6 VDD A1N hnet15 VDD LPPFET W=0.4U L=0.12U M=1 
X7 hnet15 A0N net13 VDD LPPFET W=0.4U L=0.12U M=1 
.ENDS AOI2BB1X1TS 

**** 
*.SUBCKT AOI2BB1X2TS Y A0N A1N B0 
.SUBCKT AOI2BB1X2TS Y A0N A1N B0 VSS VDD
X0 Y B0 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X1 Y net13 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X2 VDD B0 hnet10 VDD LPPFET W=0.8U L=0.12U M=1 
X3 hnet10 net13 Y VDD LPPFET W=0.8U L=0.12U M=1 
X4 VDD B0 hnet8 VDD LPPFET W=0.8U L=0.12U M=1 
X5 hnet8 net13 Y VDD LPPFET W=0.8U L=0.12U M=1 
X6 net13 A1N VSS VSS LPNFET W=0.44U L=0.12U M=1 
X7 net13 A0N VSS VSS LPNFET W=0.44U L=0.12U M=1 
X8 VDD A1N hnet16 VDD LPPFET W=0.8U L=0.12U M=1 
X9 hnet16 A0N net13 VDD LPPFET W=0.8U L=0.12U M=1 
.ENDS AOI2BB1X2TS 

**** 
*.SUBCKT AOI2BB1X4TS Y A0N A1N B0 
.SUBCKT AOI2BB1X4TS Y A0N A1N B0 VSS VDD
X0 Y B0 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X1 Y net13 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X10 VDD A1N hnet18 VDD LPPFET W=0.8U L=0.12U M=1 
X11 hnet18 A0N net13 VDD LPPFET W=0.8U L=0.12U M=1 
X12 VDD A1N hnet16 VDD LPPFET W=0.8U L=0.12U M=1 
X13 hnet16 A0N net13 VDD LPPFET W=0.8U L=0.12U M=1 
X2 VDD B0 hnet10 VDD LPPFET W=1.12U L=0.12U M=1 
X3 hnet10 net13 Y VDD LPPFET W=1.12U L=0.12U M=1 
X4 VDD B0 hnet8 VDD LPPFET W=1.12U L=0.12U M=1 
X5 hnet8 net13 Y VDD LPPFET W=1.12U L=0.12U M=1 
X6 VDD B0 hnet12 VDD LPPFET W=1.12U L=0.12U M=1 
X7 hnet12 net13 Y VDD LPPFET W=1.12U L=0.12U M=1 
X8 net13 A1N VSS VSS LPNFET W=0.78U L=0.12U M=1 
X9 net13 A0N VSS VSS LPNFET W=0.78U L=0.12U M=1 
.ENDS AOI2BB1X4TS 

**** 
*.SUBCKT AOI2BB1XLTS Y A0N A1N B0 
.SUBCKT AOI2BB1XLTS Y A0N A1N B0 VSS VDD
X0 Y B0 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X1 Y net13 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X2 VDD B0 hnet9 VDD LPPFET W=0.44U L=0.12U M=1 
X3 hnet9 net13 Y VDD LPPFET W=0.44U L=0.12U M=1 
X4 net13 A1N VSS VSS LPNFET W=0.2U L=0.12U M=1 
X5 net13 A0N VSS VSS LPNFET W=0.2U L=0.12U M=1 
X6 VDD A1N hnet15 VDD LPPFET W=0.3U L=0.12U M=1 
X7 hnet15 A0N net13 VDD LPPFET W=0.3U L=0.12U M=1 
.ENDS AOI2BB1XLTS 

**** 
*.SUBCKT AOI2BB2X1TS Y A0N A1N B0 B1 
.SUBCKT AOI2BB2X1TS Y A0N A1N B0 B1 VSS VDD
X0 hnet15 B1 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X1 Y B0 hnet15 VSS LPNFET W=0.6U L=0.12U M=1 
X2 nmin1 A1N VSS VSS LPNFET W=0.22U L=0.12U M=1 
X3 nmin1 A0N VSS VSS LPNFET W=0.22U L=0.12U M=1 
X4 VDD A1N hnet17 VDD LPPFET W=0.4U L=0.12U M=1 
X5 hnet17 A0N nmin1 VDD LPPFET W=0.4U L=0.12U M=1 
X6 Y nmin1 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X7 Y nmin1 net41 VDD LPPFET W=0.84U L=0.12U M=1 
X8 net41 B0 VDD VDD LPPFET W=0.84U L=0.12U M=1 
X9 net41 B1 VDD VDD LPPFET W=0.72U L=0.12U M=1 
.ENDS AOI2BB2X1TS 

**** 
*.SUBCKT AOI2BB2X2TS Y A0N A1N B0 B1 
.SUBCKT AOI2BB2X2TS Y A0N A1N B0 B1 VSS VDD
X0 hnet16 B1 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X1 Y B0 hnet16 VSS LPNFET W=0.6U L=0.12U M=1 
X10 net41 B0 VDD VDD LPPFET W=1.68U L=0.12U M=1 
X11 net41 B1 VDD VDD LPPFET W=1.68U L=0.12U M=1 
X2 hnet12 B1 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X3 Y B0 hnet12 VSS LPNFET W=0.6U L=0.12U M=1 
X4 nmin1 A1N VSS VSS LPNFET W=0.44U L=0.12U M=1 
X5 nmin1 A0N VSS VSS LPNFET W=0.44U L=0.12U M=1 
X6 VDD A1N hnet18 VDD LPPFET W=0.8U L=0.12U M=1 
X7 hnet18 A0N nmin1 VDD LPPFET W=0.8U L=0.12U M=1 
X8 Y nmin1 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X9 Y nmin1 net41 VDD LPPFET W=1.68U L=0.12U M=1 
.ENDS AOI2BB2X2TS 

**** 
*.SUBCKT AOI2BB2X4TS Y A0N A1N B0 B1 
.SUBCKT AOI2BB2X4TS Y A0N A1N B0 B1 VSS VDD
X0 hnet17 B1 VSS VSS LPNFET W=0.82U L=0.12U M=1 
X1 Y B0 hnet17 VSS LPNFET W=0.82U L=0.12U M=1 
X10 VDD A1N hnet18 VDD LPPFET W=0.8U L=0.12U M=1 
X11 hnet18 A0N nmin1 VDD LPPFET W=0.8U L=0.12U M=1 
X12 Y nmin1 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X13 Y nmin1 net41 VDD LPPFET W=3.36U L=0.12U M=1 
X14 net41 B0 VDD VDD LPPFET W=3.36U L=0.12U M=1 
X15 net41 B1 VDD VDD LPPFET W=3.36U L=0.12U M=1 
X2 hnet12 B1 VSS VSS LPNFET W=0.82U L=0.12U M=1 
X3 Y B0 hnet12 VSS LPNFET W=0.82U L=0.12U M=1 
X4 hnet16 B1 VSS VSS LPNFET W=0.82U L=0.12U M=1 
X5 Y B0 hnet16 VSS LPNFET W=0.82U L=0.12U M=1 
X6 nmin1 A1N VSS VSS LPNFET W=0.86U L=0.12U M=1 
X7 nmin1 A0N VSS VSS LPNFET W=0.86U L=0.12U M=1 
X8 VDD A1N hnet20 VDD LPPFET W=0.8U L=0.12U M=1 
X9 hnet20 A0N nmin1 VDD LPPFET W=0.8U L=0.12U M=1 
.ENDS AOI2BB2X4TS 

**** 
*.SUBCKT AOI2BB2XLTS Y A0N A1N B0 B1 
.SUBCKT AOI2BB2XLTS Y A0N A1N B0 B1 VSS VDD
X0 hnet15 B1 VSS VSS LPNFET W=0.4U L=0.12U M=1 
X1 Y B0 hnet15 VSS LPNFET W=0.4U L=0.12U M=1 
X2 nmin1 A1N VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 nmin1 A0N VSS VSS LPNFET W=0.2U L=0.12U M=1 
X4 VDD A1N hnet17 VDD LPPFET W=0.3U L=0.12U M=1 
X5 hnet17 A0N nmin1 VDD LPPFET W=0.3U L=0.12U M=1 
X6 Y nmin1 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X7 Y nmin1 net41 VDD LPPFET W=0.44U L=0.12U M=1 
X8 net41 B0 VDD VDD LPPFET W=0.44U L=0.12U M=1 
X9 net41 B1 VDD VDD LPPFET W=0.44U L=0.12U M=1 
.ENDS AOI2BB2XLTS 

**** 
*.SUBCKT AOI31X1TS Y A0 A1 A2 B0 
.SUBCKT AOI31X1TS Y A0 A1 A2 B0 VSS VDD
X0 hnet16 A2 VSS VSS LPNFET W=0.66U L=0.12U M=1 
X1 hnet11 A1 hnet16 VSS LPNFET W=0.66U L=0.12U M=1 
X2 Y A0 hnet11 VSS LPNFET W=0.66U L=0.12U M=1 
X3 net23 A0 VDD VDD LPPFET W=0.84U L=0.12U M=1 
X4 Y B0 net23 VDD LPPFET W=0.84U L=0.12U M=1 
X5 net23 A2 VDD VDD LPPFET W=0.84U L=0.12U M=1 
X6 net23 A1 VDD VDD LPPFET W=0.84U L=0.12U M=1 
X7 Y B0 VSS VSS LPNFET W=0.46U L=0.12U M=1 
.ENDS AOI31X1TS 

**** 
*.SUBCKT AOI31X2TS Y A0 A1 A2 B0 
.SUBCKT AOI31X2TS Y A0 A1 A2 B0 VSS VDD
X0 hnet17 A2 VSS VSS LPNFET W=0.72U L=0.12U M=1 
X1 hnet11 A1 hnet17 VSS LPNFET W=0.72U L=0.12U M=1 
X10 Y B0 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X2 Y A0 hnet11 VSS LPNFET W=0.72U L=0.12U M=1 
X3 hnet18 A2 VSS VSS LPNFET W=0.72U L=0.12U M=1 
X4 hnet13 A1 hnet18 VSS LPNFET W=0.72U L=0.12U M=1 
X5 Y A0 hnet13 VSS LPNFET W=0.72U L=0.12U M=1 
X6 net23 A0 VDD VDD LPPFET W=1.68U L=0.12U M=1 
X7 Y B0 net23 VDD LPPFET W=1.68U L=0.12U M=1 
X8 net23 A2 VDD VDD LPPFET W=1.68U L=0.12U M=1 
X9 net23 A1 VDD VDD LPPFET W=1.68U L=0.12U M=1 
.ENDS AOI31X2TS 

**** 
*.SUBCKT AOI31X4TS Y A0 A1 A2 B0 
.SUBCKT AOI31X4TS Y A0 A1 A2 B0 VSS VDD
X0 VDD net22 net18 VDD LPPFET W=1.02U L=0.12U M=1 
X1 net18 net22 VSS VSS LPNFET W=0.74U L=0.12U M=1 
X10 net28 A1 VDD VDD LPPFET W=0.54U L=0.12U M=1 
X11 net22 B0 VSS VSS LPNFET W=0.3U L=0.12U M=1 
X2 VDD net18 Y VDD LPPFET W=2.56U L=0.12U M=1 
X3 Y net18 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X4 hnet22 A2 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X5 hnet17 A1 hnet22 VSS LPNFET W=0.46U L=0.12U M=1 
X6 net22 A0 hnet17 VSS LPNFET W=0.46U L=0.12U M=1 
X7 net28 A0 VDD VDD LPPFET W=0.54U L=0.12U M=1 
X8 net22 B0 net28 VDD LPPFET W=0.54U L=0.12U M=1 
X9 net28 A2 VDD VDD LPPFET W=0.54U L=0.12U M=1 
.ENDS AOI31X4TS 

**** 
*.SUBCKT AOI31XLTS Y A0 A1 A2 B0 
.SUBCKT AOI31XLTS Y A0 A1 A2 B0 VSS VDD
X0 hnet16 A2 VSS VSS LPNFET W=0.48U L=0.12U M=1 
X1 hnet11 A1 hnet16 VSS LPNFET W=0.48U L=0.12U M=1 
X2 Y A0 hnet11 VSS LPNFET W=0.48U L=0.12U M=1 
X3 net23 A0 VDD VDD LPPFET W=0.44U L=0.12U M=1 
X4 Y B0 net23 VDD LPPFET W=0.44U L=0.12U M=1 
X5 net23 A2 VDD VDD LPPFET W=0.44U L=0.12U M=1 
X6 net23 A1 VDD VDD LPPFET W=0.44U L=0.12U M=1 
X7 Y B0 VSS VSS LPNFET W=0.24U L=0.12U M=1 
.ENDS AOI31XLTS 

**** 
*.SUBCKT AOI32X1TS Y A0 A1 A2 B0 B1 
.SUBCKT AOI32X1TS Y A0 A1 A2 B0 B1 VSS VDD
X0 hnet17 A2 VSS VSS LPNFET W=0.72U L=0.12U M=1 
X1 hnet11 A1 hnet17 VSS LPNFET W=0.72U L=0.12U M=1 
X2 Y A0 hnet11 VSS LPNFET W=0.72U L=0.12U M=1 
X3 hnet21 B1 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X4 Y B0 hnet21 VSS LPNFET W=0.6U L=0.12U M=1 
X5 net37 A0 VDD VDD LPPFET W=0.84U L=0.12U M=1 
X6 net37 A1 VDD VDD LPPFET W=0.84U L=0.12U M=1 
X7 Y B0 net37 VDD LPPFET W=0.84U L=0.12U M=1 
X8 net37 A2 VDD VDD LPPFET W=0.84U L=0.12U M=1 
X9 Y B1 net37 VDD LPPFET W=0.84U L=0.12U M=1 
.ENDS AOI32X1TS 

**** 
*.SUBCKT AOI32X2TS Y A0 A1 A2 B0 B1 
.SUBCKT AOI32X2TS Y A0 A1 A2 B0 B1 VSS VDD
X0 hnet18 A2 VSS VSS LPNFET W=0.7U L=0.12U M=1 
X1 hnet11 A1 hnet18 VSS LPNFET W=0.7U L=0.12U M=1 
X10 net37 A0 VDD VDD LPPFET W=1.68U L=0.12U M=1 
X11 net37 A1 VDD VDD LPPFET W=1.68U L=0.12U M=1 
X12 Y B0 net37 VDD LPPFET W=1.52U L=0.12U M=1 
X13 net37 A2 VDD VDD LPPFET W=1.68U L=0.12U M=1 
X14 Y B1 net37 VDD LPPFET W=1.68U L=0.12U M=1 
X2 Y A0 hnet11 VSS LPNFET W=0.7U L=0.12U M=1 
X3 hnet19 A2 VSS VSS LPNFET W=0.7U L=0.12U M=1 
X4 hnet14 A1 hnet19 VSS LPNFET W=0.7U L=0.12U M=1 
X5 Y A0 hnet14 VSS LPNFET W=0.7U L=0.12U M=1 
X6 hnet24 B1 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X7 Y B0 hnet24 VSS LPNFET W=0.6U L=0.12U M=1 
X8 hnet20 B1 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X9 Y B0 hnet20 VSS LPNFET W=0.6U L=0.12U M=1 
.ENDS AOI32X2TS 

**** 
*.SUBCKT AOI32X4TS Y A0 A1 A2 B0 B1 
.SUBCKT AOI32X4TS Y A0 A1 A2 B0 B1 VSS VDD
X0 VDD net24 net20 VDD LPPFET W=1.02U L=0.12U M=1 
X1 net20 net24 VSS VSS LPNFET W=0.74U L=0.12U M=1 
X10 net42 A1 VDD VDD LPPFET W=0.54U L=0.12U M=1 
X11 net24 B0 net42 VDD LPPFET W=0.54U L=0.12U M=1 
X12 net42 A2 VDD VDD LPPFET W=0.54U L=0.12U M=1 
X13 net24 B1 net42 VDD LPPFET W=0.54U L=0.12U M=1 
X2 VDD net20 Y VDD LPPFET W=2.56U L=0.12U M=1 
X3 Y net20 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X4 hnet24 A2 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X5 hnet19 A1 hnet24 VSS LPNFET W=0.46U L=0.12U M=1 
X6 net24 A0 hnet19 VSS LPNFET W=0.46U L=0.12U M=1 
X7 hnet28 B1 VSS VSS LPNFET W=0.38U L=0.12U M=1 
X8 net24 B0 hnet28 VSS LPNFET W=0.38U L=0.12U M=1 
X9 net42 A0 VDD VDD LPPFET W=0.54U L=0.12U M=1 
.ENDS AOI32X4TS 

**** 
*.SUBCKT AOI32XLTS Y A0 A1 A2 B0 B1 
.SUBCKT AOI32XLTS Y A0 A1 A2 B0 B1 VSS VDD
X0 hnet17 A2 VSS VSS LPNFET W=0.48U L=0.12U M=1 
X1 hnet11 A1 hnet17 VSS LPNFET W=0.48U L=0.12U M=1 
X2 Y A0 hnet11 VSS LPNFET W=0.48U L=0.12U M=1 
X3 hnet21 B1 VSS VSS LPNFET W=0.4U L=0.12U M=1 
X4 Y B0 hnet21 VSS LPNFET W=0.4U L=0.12U M=1 
X5 net37 A0 VDD VDD LPPFET W=0.44U L=0.12U M=1 
X6 net37 A1 VDD VDD LPPFET W=0.44U L=0.12U M=1 
X7 Y B0 net37 VDD LPPFET W=0.44U L=0.12U M=1 
X8 net37 A2 VDD VDD LPPFET W=0.44U L=0.12U M=1 
X9 Y B1 net37 VDD LPPFET W=0.44U L=0.12U M=1 
.ENDS AOI32XLTS 

**** 
*.SUBCKT AOI33X1TS Y A0 A1 A2 B0 B1 B2 
.SUBCKT AOI33X1TS Y A0 A1 A2 B0 B1 B2 VSS VDD
X0 hnet18 B2 VSS VSS LPNFET W=0.72U L=0.12U M=1 
X1 hnet12 B1 hnet18 VSS LPNFET W=0.72U L=0.12U M=1 
X10 net46 B2 VDD VDD LPPFET W=0.84U L=0.12U M=1 
X11 Y A2 net46 VDD LPPFET W=0.84U L=0.12U M=1 
X2 Y B0 hnet12 VSS LPNFET W=0.72U L=0.12U M=1 
X3 hnet25 A2 VSS VSS LPNFET W=0.72U L=0.12U M=1 
X4 hnet19 A1 hnet25 VSS LPNFET W=0.72U L=0.12U M=1 
X5 Y A0 hnet19 VSS LPNFET W=0.72U L=0.12U M=1 
X6 net46 B0 VDD VDD LPPFET W=0.84U L=0.12U M=1 
X7 Y A0 net46 VDD LPPFET W=0.84U L=0.12U M=1 
X8 net46 B1 VDD VDD LPPFET W=0.84U L=0.12U M=1 
X9 Y A1 net46 VDD LPPFET W=0.84U L=0.12U M=1 
.ENDS AOI33X1TS 

**** 
*.SUBCKT AOI33X2TS Y A0 A1 A2 B0 B1 B2 
.SUBCKT AOI33X2TS Y A0 A1 A2 B0 B1 B2 VSS VDD
X0 hnet19 B2 VSS VSS LPNFET W=0.72U L=0.12U M=1 
X1 hnet12 B1 hnet19 VSS LPNFET W=0.72U L=0.12U M=1 
X10 hnet24 A1 hnet29 VSS LPNFET W=0.72U L=0.12U M=1 
X11 Y A0 hnet24 VSS LPNFET W=0.72U L=0.12U M=1 
X12 net46 B0 VDD VDD LPPFET W=1.68U L=0.12U M=1 
X13 Y A0 net46 VDD LPPFET W=1.68U L=0.12U M=1 
X14 net46 B1 VDD VDD LPPFET W=1.68U L=0.12U M=1 
X15 Y A1 net46 VDD LPPFET W=1.68U L=0.12U M=1 
X16 net46 B2 VDD VDD LPPFET W=1.68U L=0.12U M=1 
X17 Y A2 net46 VDD LPPFET W=1.68U L=0.12U M=1 
X2 Y B0 hnet12 VSS LPNFET W=0.72U L=0.12U M=1 
X3 hnet20 B2 VSS VSS LPNFET W=0.72U L=0.12U M=1 
X4 hnet15 B1 hnet20 VSS LPNFET W=0.72U L=0.12U M=1 
X5 Y B0 hnet15 VSS LPNFET W=0.72U L=0.12U M=1 
X6 hnet28 A2 VSS VSS LPNFET W=0.72U L=0.12U M=1 
X7 hnet21 A1 hnet28 VSS LPNFET W=0.72U L=0.12U M=1 
X8 Y A0 hnet21 VSS LPNFET W=0.72U L=0.12U M=1 
X9 hnet29 A2 VSS VSS LPNFET W=0.72U L=0.12U M=1 
.ENDS AOI33X2TS 

**** 
*.SUBCKT AOI33X4TS Y A0 A1 A2 B0 B1 B2 
.SUBCKT AOI33X4TS Y A0 A1 A2 B0 B1 B2 VSS VDD
X0 VDD net27 Y VDD LPPFET W=2.56U L=0.12U M=1 
X1 Y net27 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X10 net51 B0 VDD VDD LPPFET W=0.54U L=0.12U M=1 
X11 net29 A0 net51 VDD LPPFET W=0.54U L=0.12U M=1 
X12 net51 B1 VDD VDD LPPFET W=0.54U L=0.12U M=1 
X13 net29 A1 net51 VDD LPPFET W=0.54U L=0.12U M=1 
X14 net51 B2 VDD VDD LPPFET W=0.54U L=0.12U M=1 
X15 net29 A2 net51 VDD LPPFET W=0.54U L=0.12U M=1 
X2 VDD net29 net27 VDD LPPFET W=1.02U L=0.12U M=1 
X3 net27 net29 VSS VSS LPNFET W=0.74U L=0.12U M=1 
X4 hnet25 B2 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X5 hnet20 B1 hnet25 VSS LPNFET W=0.46U L=0.12U M=1 
X6 net29 B0 hnet20 VSS LPNFET W=0.46U L=0.12U M=1 
X7 hnet31 A2 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X8 hnet26 A1 hnet31 VSS LPNFET W=0.46U L=0.12U M=1 
X9 net29 A0 hnet26 VSS LPNFET W=0.46U L=0.12U M=1 
.ENDS AOI33X4TS 

**** 
*.SUBCKT AOI33XLTS Y A0 A1 A2 B0 B1 B2 
.SUBCKT AOI33XLTS Y A0 A1 A2 B0 B1 B2 VSS VDD
X0 hnet18 B2 VSS VSS LPNFET W=0.48U L=0.12U M=1 
X1 hnet12 B1 hnet18 VSS LPNFET W=0.48U L=0.12U M=1 
X10 net46 B2 VDD VDD LPPFET W=0.44U L=0.12U M=1 
X11 Y A2 net46 VDD LPPFET W=0.44U L=0.12U M=1 
X2 Y B0 hnet12 VSS LPNFET W=0.48U L=0.12U M=1 
X3 hnet25 A2 VSS VSS LPNFET W=0.48U L=0.12U M=1 
X4 hnet19 A1 hnet25 VSS LPNFET W=0.48U L=0.12U M=1 
X5 Y A0 hnet19 VSS LPNFET W=0.48U L=0.12U M=1 
X6 net46 B0 VDD VDD LPPFET W=0.44U L=0.12U M=1 
X7 Y A0 net46 VDD LPPFET W=0.44U L=0.12U M=1 
X8 net46 B1 VDD VDD LPPFET W=0.44U L=0.12U M=1 
X9 Y A1 net46 VDD LPPFET W=0.44U L=0.12U M=1 
.ENDS AOI33XLTS 

**** 
*.SUBCKT BENCX1TS A S X2 M0 M1 M2 
.SUBCKT BENCX1TS A S X2 M0 M1 M2 VSS VDD
X0 VDD nm1 hnet26 VDD LPPFET W=0.56U L=0.12U M=1 
X1 hnet26 nm0 net60 VDD LPPFET W=0.56U L=0.12U M=1 
X10 net78 nm1 VSS VSS LPNFET W=0.34U L=0.12U M=1 
X11 net63 nm2 net87 VSS LPNFET W=0.34U L=0.12U M=1 
X12 net87 M0 VSS VSS LPNFET W=0.34U L=0.12U M=1 
X13 net87 M1 VSS VSS LPNFET W=0.34U L=0.12U M=1 
X14 net93 nm1 nm0 VSS LPNFET W=0.34U L=0.12U M=1 
X15 net93 M1 net106 VSS LPNFET W=0.34U L=0.12U M=1 
X16 VDD net102 S VDD LPPFET W=2.6U L=0.12U M=1 
X17 S net102 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X18 VDD net104 A VDD LPPFET W=2.6U L=0.12U M=1 
X19 A net104 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X2 VDD M1 hnet30 VDD LPPFET W=0.56U L=0.12U M=1 
X20 VDD net112 X2 VDD LPPFET W=2.6U L=0.12U M=1 
X21 X2 net112 VSS VSS LPNFET W=1.66U L=0.12U M=1 
X22 VDD M2 nm2 VDD LPPFET W=0.28U L=0.12U M=1 
X23 nm2 M2 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X24 VDD net60 net102 VDD LPPFET W=0.78U L=0.12U M=1 
X25 net102 net60 VSS VSS LPNFET W=0.56U L=0.12U M=1 
X26 VDD net63 net104 VDD LPPFET W=0.78U L=0.12U M=1 
X27 net104 net63 VSS VSS LPNFET W=0.56U L=0.12U M=1 
X28 VDD nm0 net106 VDD LPPFET W=0.48U L=0.12U M=1 
X29 net106 nm0 VSS VSS LPNFET W=0.34U L=0.12U M=1 
X3 hnet30 M0 net63 VDD LPPFET W=0.56U L=0.12U M=1 
X30 VDD M1 nm1 VDD LPPFET W=0.3U L=0.12U M=1 
X31 nm1 M1 VSS VSS LPNFET W=0.22U L=0.12U M=1 
X32 VDD M0 nm0 VDD LPPFET W=0.78U L=0.12U M=1 
X33 nm0 M0 VSS VSS LPNFET W=0.56U L=0.12U M=1 
X34 VDD net93 net112 VDD LPPFET W=0.78U L=0.12U M=1 
X35 net112 net93 VSS VSS LPNFET W=0.56U L=0.12U M=1 
X4 net60 M2 VDD VDD LPPFET W=0.28U L=0.12U M=1 
X5 net63 nm2 VDD VDD LPPFET W=0.28U L=0.12U M=1 
X6 net93 M1 nm0 VDD LPPFET W=0.48U L=0.12U M=1 
X7 net93 nm1 net106 VDD LPPFET W=0.48U L=0.12U M=1 
X8 net60 M2 net78 VSS LPNFET W=0.3U L=0.12U M=1 
X9 net78 nm0 VSS VSS LPNFET W=0.34U L=0.12U M=1 
.ENDS BENCX1TS 

**** 
*.SUBCKT BENCX2TS A S X2 M0 M1 M2 
.SUBCKT BENCX2TS A S X2 M0 M1 M2 VSS VDD
X0 VDD nm1 hnet26 VDD LPPFET W=1U L=0.12U M=1 
X1 hnet26 nm0 net60 VDD LPPFET W=1U L=0.12U M=1 
X10 net78 nm1 VSS VSS LPNFET W=0.68U L=0.12U M=1 
X11 net63 nm2 net87 VSS LPNFET W=0.68U L=0.12U M=1 
X12 net87 M0 VSS VSS LPNFET W=0.68U L=0.12U M=1 
X13 net87 M1 VSS VSS LPNFET W=0.68U L=0.12U M=1 
X14 net93 nm1 nm0 VSS LPNFET W=0.66U L=0.12U M=1 
X15 net93 M1 net106 VSS LPNFET W=0.66U L=0.12U M=1 
X16 VDD net102 S VDD LPPFET W=5.2U L=0.12U M=1 
X17 S net102 VSS VSS LPNFET W=3.68U L=0.12U M=1 
X18 VDD net104 A VDD LPPFET W=5.2U L=0.12U M=1 
X19 A net104 VSS VSS LPNFET W=3.68U L=0.12U M=1 
X2 VDD M1 hnet30 VDD LPPFET W=1U L=0.12U M=1 
X20 VDD net112 X2 VDD LPPFET W=5.2U L=0.12U M=1 
X21 X2 net112 VSS VSS LPNFET W=3.24U L=0.12U M=1 
X22 VDD M2 nm2 VDD LPPFET W=0.28U L=0.12U M=1 
X23 nm2 M2 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X24 VDD net60 net102 VDD LPPFET W=1.56U L=0.12U M=1 
X25 net102 net60 VSS VSS LPNFET W=1.12U L=0.12U M=1 
X26 VDD net63 net104 VDD LPPFET W=1.56U L=0.12U M=1 
X27 net104 net63 VSS VSS LPNFET W=1.12U L=0.12U M=1 
X28 VDD nm0 net106 VDD LPPFET W=0.94U L=0.12U M=1 
X29 net106 nm0 VSS VSS LPNFET W=0.68U L=0.12U M=1 
X3 hnet30 M0 net63 VDD LPPFET W=1U L=0.12U M=1 
X30 VDD M1 nm1 VDD LPPFET W=0.58U L=0.12U M=1 
X31 nm1 M1 VSS VSS LPNFET W=0.42U L=0.12U M=1 
X32 VDD M0 nm0 VDD LPPFET W=1.5U L=0.12U M=1 
X33 nm0 M0 VSS VSS LPNFET W=1.08U L=0.12U M=1 
X34 VDD net93 net112 VDD LPPFET W=1.56U L=0.12U M=1 
X35 net112 net93 VSS VSS LPNFET W=1.08U L=0.12U M=1 
X4 net60 M2 VDD VDD LPPFET W=0.5U L=0.12U M=1 
X5 net63 nm2 VDD VDD LPPFET W=0.5U L=0.12U M=1 
X6 net93 M1 nm0 VDD LPPFET W=0.94U L=0.12U M=1 
X7 net93 nm1 net106 VDD LPPFET W=0.94U L=0.12U M=1 
X8 net60 M2 net78 VSS LPNFET W=0.68U L=0.12U M=1 
X9 net78 nm0 VSS VSS LPNFET W=0.68U L=0.12U M=1 
.ENDS BENCX2TS 

**** 
*.SUBCKT BENCX4TS A S X2 M0 M1 M2 
.SUBCKT BENCX4TS A S X2 M0 M1 M2 VSS VDD
X0 VDD nm1 hnet27 VDD LPPFET W=1U L=0.12U M=1 
X1 hnet27 nm0 net60 VDD LPPFET W=1U L=0.12U M=1 
X10 net93 M1 nm0 VDD LPPFET W=1.84U L=0.12U M=1 
X11 net93 nm1 net106 VDD LPPFET W=1.84U L=0.12U M=1 
X12 net60 M2 net78 VSS LPNFET W=1.44U L=0.12U M=1 
X13 net78 nm0 VSS VSS LPNFET W=1.32U L=0.12U M=1 
X14 net78 nm1 VSS VSS LPNFET W=1.32U L=0.12U M=1 
X15 net63 nm2 net87 VSS LPNFET W=1.32U L=0.12U M=1 
X16 net87 M0 VSS VSS LPNFET W=1.32U L=0.12U M=1 
X17 net87 M1 VSS VSS LPNFET W=1.32U L=0.12U M=1 
X18 net93 nm1 nm0 VSS LPNFET W=1.2U L=0.12U M=1 
X19 net93 M1 net106 VSS LPNFET W=1.32U L=0.12U M=1 
X2 VDD nm1 hnet24 VDD LPPFET W=1U L=0.12U M=1 
X20 VDD net102 S VDD LPPFET W=10.4U L=0.12U M=1 
X21 S net102 VSS VSS LPNFET W=7.1U L=0.12U M=1 
X22 VDD net104 A VDD LPPFET W=10.4U L=0.12U M=1 
X23 A net104 VSS VSS LPNFET W=7.36U L=0.12U M=1 
X24 VDD net112 X2 VDD LPPFET W=10.4U L=0.12U M=1 
X25 X2 net112 VSS VSS LPNFET W=6.96U L=0.12U M=1 
X26 VDD M2 nm2 VDD LPPFET W=0.38U L=0.12U M=1 
X27 nm2 M2 VSS VSS LPNFET W=0.28U L=0.12U M=1 
X28 VDD net60 net102 VDD LPPFET W=3.08U L=0.12U M=1 
X29 net102 net60 VSS VSS LPNFET W=2.24U L=0.12U M=1 
X3 hnet24 nm0 net60 VDD LPPFET W=1U L=0.12U M=1 
X30 VDD net63 net104 VDD LPPFET W=3.08U L=0.12U M=1 
X31 net104 net63 VSS VSS LPNFET W=2.24U L=0.12U M=1 
X32 VDD nm0 net106 VDD LPPFET W=1.84U L=0.12U M=1 
X33 net106 nm0 VSS VSS LPNFET W=1.32U L=0.12U M=1 
X34 VDD M1 nm1 VDD LPPFET W=1.12U L=0.12U M=1 
X35 nm1 M1 VSS VSS LPNFET W=0.8U L=0.12U M=1 
X36 VDD M0 nm0 VDD LPPFET W=2.98U L=0.12U M=1 
X37 nm0 M0 VSS VSS LPNFET W=2.1U L=0.12U M=1 
X38 VDD net93 net112 VDD LPPFET W=3.08U L=0.12U M=1 
X39 net112 net93 VSS VSS LPNFET W=2.22U L=0.12U M=1 
X4 VDD M1 hnet32 VDD LPPFET W=1U L=0.12U M=1 
X5 hnet32 M0 net63 VDD LPPFET W=1U L=0.12U M=1 
X6 VDD M1 hnet29 VDD LPPFET W=1U L=0.12U M=1 
X7 hnet29 M0 net63 VDD LPPFET W=1U L=0.12U M=1 
X8 net60 M2 VDD VDD LPPFET W=1U L=0.12U M=1 
X9 net63 nm2 VDD VDD LPPFET W=1U L=0.12U M=1 
.ENDS BENCX4TS 

**** 
*.SUBCKT BMXIX2TS PPN A M0 M1 S X2 
.SUBCKT BMXIX2TS PPN A M0 M1 S X2 VSS VDD
X0 VDD M1 nma1 VDD LPPFET W=0.3U L=0.12U M=1 
X1 nma1 M1 VSS VSS LPNFET W=0.22U L=0.12U M=1 
X10 VDD X2 nmx2 VDD LPPFET W=0.3U L=0.12U M=1 
X11 nmx2 X2 VSS VSS LPNFET W=0.22U L=0.12U M=1 
X12 net91 M1 nmsubb VDD LPPFET W=0.76U L=0.12U M=1 
X13 net91 nma1 nmaddb VDD LPPFET W=0.76U L=0.12U M=1 
X14 net97 M0 nmsubb VDD LPPFET W=0.74U L=0.12U M=1 
X15 net97 nma0 nmaddb VDD LPPFET W=0.7U L=0.12U M=1 
X16 net103 X2 net91 VDD LPPFET W=0.76U L=0.12U M=1 
X17 net103 nmx2 net97 VDD LPPFET W=0.76U L=0.12U M=1 
X18 net91 nma1 nmsubb VSS LPNFET W=0.56U L=0.12U M=1 
X19 net91 M1 nmaddb VSS LPNFET W=0.56U L=0.12U M=1 
X2 VDD M0 nma0 VDD LPPFET W=0.3U L=0.12U M=1 
X20 net97 nma0 nmsubb VSS LPNFET W=0.56U L=0.12U M=1 
X21 net97 M0 nmaddb VSS LPNFET W=0.56U L=0.12U M=1 
X22 net103 nmx2 net91 VSS LPNFET W=0.56U L=0.12U M=1 
X23 net103 X2 net97 VSS LPNFET W=0.56U L=0.12U M=1 
X3 nma0 M0 VSS VSS LPNFET W=0.22U L=0.12U M=1 
X4 VDD A nmaddb VDD LPPFET W=1.54U L=0.12U M=1 
X5 nmaddb A VSS VSS LPNFET W=1.1U L=0.12U M=1 
X6 VDD S nmsubb VDD LPPFET W=1.54U L=0.12U M=1 
X7 nmsubb S VSS VSS LPNFET W=1.1U L=0.12U M=1 
X8 VDD net103 PPN VDD LPPFET W=1.28U L=0.12U M=1 
X9 PPN net103 VSS VSS LPNFET W=0.92U L=0.12U M=1 
.ENDS BMXIX2TS 

**** 
*.SUBCKT BMXIX4TS PPN A M0 M1 S X2 
.SUBCKT BMXIX4TS PPN A M0 M1 S X2 VSS VDD
X0 VDD M1 nma1 VDD LPPFET W=0.62U L=0.12U M=1 
X1 nma1 M1 VSS VSS LPNFET W=0.44U L=0.12U M=1 
X10 VDD X2 nmx2 VDD LPPFET W=0.62U L=0.12U M=1 
X11 nmx2 X2 VSS VSS LPNFET W=0.44U L=0.12U M=1 
X12 net91 M1 nmsubb VDD LPPFET W=1.52U L=0.12U M=1 
X13 net91 nma1 nmaddb VDD LPPFET W=1.52U L=0.12U M=1 
X14 net97 M0 nmsubb VDD LPPFET W=1.52U L=0.12U M=1 
X15 net97 nma0 nmaddb VDD LPPFET W=1.52U L=0.12U M=1 
X16 net103 X2 net91 VDD LPPFET W=1.52U L=0.12U M=1 
X17 net103 nmx2 net97 VDD LPPFET W=1.52U L=0.12U M=1 
X18 net91 nma1 nmsubb VSS LPNFET W=1.1U L=0.12U M=1 
X19 net91 M1 nmaddb VSS LPNFET W=1.1U L=0.12U M=1 
X2 VDD M0 nma0 VDD LPPFET W=0.62U L=0.12U M=1 
X20 net97 nma0 nmsubb VSS LPNFET W=1.1U L=0.12U M=1 
X21 net97 M0 nmaddb VSS LPNFET W=1.1U L=0.12U M=1 
X22 net103 nmx2 net91 VSS LPNFET W=1.1U L=0.12U M=1 
X23 net103 X2 net97 VSS LPNFET W=1.1U L=0.12U M=1 
X3 nma0 M0 VSS VSS LPNFET W=0.44U L=0.12U M=1 
X4 VDD A nmaddb VDD LPPFET W=3.06U L=0.12U M=1 
X5 nmaddb A VSS VSS LPNFET W=2.22U L=0.12U M=1 
X6 VDD S nmsubb VDD LPPFET W=3.06U L=0.12U M=1 
X7 nmsubb S VSS VSS LPNFET W=2.2U L=0.12U M=1 
X8 VDD net103 PPN VDD LPPFET W=2.56U L=0.12U M=1 
X9 PPN net103 VSS VSS LPNFET W=1.84U L=0.12U M=1 
.ENDS BMXIX4TS 

**** 
*.SUBCKT BMXX2TS PP A M0 M1 S X2 
.SUBCKT BMXX2TS PP A M0 M1 S X2 VSS VDD
X0 VDD net103 net58 VDD LPPFET W=1.04U L=0.12U M=1 
X1 net58 net103 VSS VSS LPNFET W=0.72U L=0.12U M=1 
X10 VDD S nmsubb VDD LPPFET W=1.64U L=0.12U M=1 
X11 nmsubb S VSS VSS LPNFET W=1.18U L=0.12U M=1 
X12 VDD net109 PP VDD LPPFET W=1.28U L=0.12U M=1 
X13 PP net109 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X14 VDD X2 nmx2 VDD LPPFET W=0.42U L=0.12U M=1 
X15 nmx2 X2 VSS VSS LPNFET W=0.3U L=0.12U M=1 
X16 net97 M1 nmsubb VDD LPPFET W=0.82U L=0.12U M=1 
X17 net97 nma1 nmaddb VDD LPPFET W=0.82U L=0.12U M=1 
X18 net103 M0 nmsubb VDD LPPFET W=0.82U L=0.12U M=1 
X19 net103 nma0 nmaddb VDD LPPFET W=0.76U L=0.12U M=1 
X2 VDD net97 net60 VDD LPPFET W=1.04U L=0.12U M=1 
X20 net109 X2 net60 VDD LPPFET W=1.04U L=0.12U M=1 
X21 net109 nmx2 net58 VDD LPPFET W=0.98U L=0.12U M=1 
X22 net97 nma1 nmsubb VSS LPNFET W=0.6U L=0.12U M=1 
X23 net97 M1 nmaddb VSS LPNFET W=0.6U L=0.12U M=1 
X24 net103 nma0 nmsubb VSS LPNFET W=0.6U L=0.12U M=1 
X25 net103 M0 nmaddb VSS LPNFET W=0.6U L=0.12U M=1 
X26 net109 nmx2 net60 VSS LPNFET W=0.72U L=0.12U M=1 
X27 net109 X2 net58 VSS LPNFET W=0.74U L=0.12U M=1 
X3 net60 net97 VSS VSS LPNFET W=0.72U L=0.12U M=1 
X4 VDD M1 nma1 VDD LPPFET W=0.34U L=0.12U M=1 
X5 nma1 M1 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X6 VDD M0 nma0 VDD LPPFET W=0.34U L=0.12U M=1 
X7 nma0 M0 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X8 VDD A nmaddb VDD LPPFET W=1.64U L=0.12U M=1 
X9 nmaddb A VSS VSS LPNFET W=1.18U L=0.12U M=1 
.ENDS BMXX2TS 

**** 
*.SUBCKT BMXX4TS PP A M0 M1 S X2 
.SUBCKT BMXX4TS PP A M0 M1 S X2 VSS VDD
X0 VDD net103 net58 VDD LPPFET W=2.06U L=0.12U M=1 
X1 net58 net103 VSS VSS LPNFET W=1.48U L=0.12U M=1 
X10 VDD S nmsubb VDD LPPFET W=3.28U L=0.12U M=1 
X11 nmsubb S VSS VSS LPNFET W=2.36U L=0.12U M=1 
X12 VDD net109 PP VDD LPPFET W=2.56U L=0.12U M=1 
X13 PP net109 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X14 VDD X2 nmx2 VDD LPPFET W=0.84U L=0.12U M=1 
X15 nmx2 X2 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X16 net97 M1 nmsubb VDD LPPFET W=1.64U L=0.12U M=1 
X17 net97 nma1 nmaddb VDD LPPFET W=1.64U L=0.12U M=1 
X18 net103 M0 nmsubb VDD LPPFET W=1.64U L=0.12U M=1 
X19 net103 nma0 nmaddb VDD LPPFET W=1.64U L=0.12U M=1 
X2 VDD net97 net60 VDD LPPFET W=2.06U L=0.12U M=1 
X20 net109 X2 net60 VDD LPPFET W=2.06U L=0.12U M=1 
X21 net109 nmx2 net58 VDD LPPFET W=1.96U L=0.12U M=1 
X22 net97 nma1 nmsubb VSS LPNFET W=1.14U L=0.12U M=1 
X23 net97 M1 nmaddb VSS LPNFET W=1.1U L=0.12U M=1 
X24 net103 nma0 nmsubb VSS LPNFET W=1.18U L=0.12U M=1 
X25 net103 M0 nmaddb VSS LPNFET W=1.14U L=0.12U M=1 
X26 net109 nmx2 net60 VSS LPNFET W=1.48U L=0.12U M=1 
X27 net109 X2 net58 VSS LPNFET W=1.48U L=0.12U M=1 
X3 net60 net97 VSS VSS LPNFET W=1.48U L=0.12U M=1 
X4 VDD M1 nma1 VDD LPPFET W=0.66U L=0.12U M=1 
X5 nma1 M1 VSS VSS LPNFET W=0.48U L=0.12U M=1 
X6 VDD M0 nma0 VDD LPPFET W=0.66U L=0.12U M=1 
X7 nma0 M0 VSS VSS LPNFET W=0.48U L=0.12U M=1 
X8 VDD A nmaddb VDD LPPFET W=3.28U L=0.12U M=1 
X9 nmaddb A VSS VSS LPNFET W=2.4U L=0.12U M=1 
.ENDS BMXX4TS 

**** 
*.SUBCKT BUFX12TS Y A 
.SUBCKT BUFX12TS Y A VSS VDD
X0 VDD nmin Y VDD LPPFET W=7.24U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=4.84U L=0.12U M=1 
X2 VDD A nmin VDD LPPFET W=2.6U L=0.12U M=1 
X3 nmin A VSS VSS LPNFET W=1.84U L=0.12U M=1 
.ENDS BUFX12TS 

**** 
*.SUBCKT BUFX16TS Y A 
.SUBCKT BUFX16TS Y A VSS VDD
X0 VDD nmin Y VDD LPPFET W=9.88U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=6.8U L=0.12U M=1 
X2 VDD A nmin VDD LPPFET W=3.9U L=0.12U M=1 
X3 nmin A VSS VSS LPNFET W=2.76U L=0.12U M=1 
.ENDS BUFX16TS 

**** 
*.SUBCKT BUFX20TS Y A 
.SUBCKT BUFX20TS Y A VSS VDD
X0 VDD nmin Y VDD LPPFET W=12.74U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=8.94U L=0.12U M=1 
X2 VDD A nmin VDD LPPFET W=5.12U L=0.12U M=1 
X3 nmin A VSS VSS LPNFET W=3.68U L=0.12U M=1 
.ENDS BUFX20TS 

**** 
*.SUBCKT BUFX2TS Y A 
.SUBCKT BUFX2TS Y A VSS VDD
X0 VDD nmin Y VDD LPPFET W=1.28U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=0.92U L=0.12U M=1 
X2 VDD A nmin VDD LPPFET W=0.5U L=0.12U M=1 
X3 nmin A VSS VSS LPNFET W=0.34U L=0.12U M=1 
.ENDS BUFX2TS 

**** 
*.SUBCKT BUFX3TS Y A 
.SUBCKT BUFX3TS Y A VSS VDD
X0 VDD nmin Y VDD LPPFET W=1.92U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=1.38U L=0.12U M=1 
X2 VDD A nmin VDD LPPFET W=0.78U L=0.12U M=1 
X3 nmin A VSS VSS LPNFET W=0.56U L=0.12U M=1 
.ENDS BUFX3TS 

**** 
*.SUBCKT BUFX4TS Y A 
.SUBCKT BUFX4TS Y A VSS VDD
X0 VDD nmin Y VDD LPPFET W=2.56U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=1.84U L=0.12U M=1 
X2 VDD A nmin VDD LPPFET W=1.02U L=0.12U M=1 
X3 nmin A VSS VSS LPNFET W=0.68U L=0.12U M=1 
.ENDS BUFX4TS 

**** 
*.SUBCKT BUFX6TS Y A 
.SUBCKT BUFX6TS Y A VSS VDD
X0 VDD nmin Y VDD LPPFET W=3.84U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=2.76U L=0.12U M=1 
X2 VDD A nmin VDD LPPFET W=1.54U L=0.12U M=1 
X3 nmin A VSS VSS LPNFET W=1.1U L=0.12U M=1 
.ENDS BUFX6TS 

**** 
*.SUBCKT BUFX8TS Y A 
.SUBCKT BUFX8TS Y A VSS VDD
X0 VDD nmin Y VDD LPPFET W=5.12U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=3.68U L=0.12U M=1 
X2 VDD A nmin VDD LPPFET W=2.06U L=0.12U M=1 
X3 nmin A VSS VSS LPNFET W=1.34U L=0.12U M=1 
.ENDS BUFX8TS 

**** 
*.SUBCKT CLKAND2X12TS Y A B 
.SUBCKT CLKAND2X12TS Y A B VSS VDD
X0 VDD net11 Y VDD LPPFET W=6.76U L=0.12U M=1 
X1 Y net11 VSS VSS LPNFET W=2.56U L=0.12U M=1 
X2 hnet15 B VSS VSS LPNFET W=0.56U L=0.12U M=1 
X3 net11 A hnet15 VSS LPNFET W=0.56U L=0.12U M=1 
X4 hnet11 B VSS VSS LPNFET W=0.56U L=0.12U M=1 
X5 net11 A hnet11 VSS LPNFET W=0.56U L=0.12U M=1 
X6 VDD B net11 VDD LPPFET W=2.94U L=0.12U M=1 
X7 VDD A net11 VDD LPPFET W=2.94U L=0.12U M=1 
.ENDS CLKAND2X12TS 

**** 
*.SUBCKT CLKAND2X2TS Y A B 
.SUBCKT CLKAND2X2TS Y A B VSS VDD
X0 VDD net11 Y VDD LPPFET W=1.3U L=0.12U M=1 
X1 Y net11 VSS VSS LPNFET W=0.48U L=0.12U M=1 
X2 hnet14 B VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 net11 A hnet14 VSS LPNFET W=0.2U L=0.12U M=1 
X4 VDD B net11 VDD LPPFET W=0.56U L=0.12U M=1 
X5 VDD A net11 VDD LPPFET W=0.56U L=0.12U M=1 
.ENDS CLKAND2X2TS 

**** 
*.SUBCKT CLKAND2X3TS Y A B 
.SUBCKT CLKAND2X3TS Y A B VSS VDD
X0 VDD net11 Y VDD LPPFET W=1.94U L=0.12U M=1 
X1 Y net11 VSS VSS LPNFET W=0.72U L=0.12U M=1 
X2 hnet14 B VSS VSS LPNFET W=0.28U L=0.12U M=1 
X3 net11 A hnet14 VSS LPNFET W=0.28U L=0.12U M=1 
X4 VDD B net11 VDD LPPFET W=0.78U L=0.12U M=1 
X5 VDD A net11 VDD LPPFET W=0.78U L=0.12U M=1 
.ENDS CLKAND2X3TS 

**** 
*.SUBCKT CLKAND2X4TS Y A B 
.SUBCKT CLKAND2X4TS Y A B VSS VDD
X0 VDD net11 Y VDD LPPFET W=2.54U L=0.12U M=1 
X1 Y net11 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X2 hnet14 B VSS VSS LPNFET W=0.36U L=0.12U M=1 
X3 net11 A hnet14 VSS LPNFET W=0.36U L=0.12U M=1 
X4 VDD B net11 VDD LPPFET W=1U L=0.12U M=1 
X5 VDD A net11 VDD LPPFET W=1U L=0.12U M=1 
.ENDS CLKAND2X4TS 

**** 
*.SUBCKT CLKAND2X6TS Y A B 
.SUBCKT CLKAND2X6TS Y A B VSS VDD
X0 VDD net11 Y VDD LPPFET W=3.02U L=0.12U M=1 
X1 Y net11 VSS VSS LPNFET W=1.12U L=0.12U M=1 
X2 hnet14 B VSS VSS LPNFET W=0.46U L=0.12U M=1 
X3 net11 A hnet14 VSS LPNFET W=0.46U L=0.12U M=1 
X4 VDD B net11 VDD LPPFET W=1.3U L=0.12U M=1 
X5 VDD A net11 VDD LPPFET W=1.3U L=0.12U M=1 
.ENDS CLKAND2X6TS 

**** 
*.SUBCKT CLKAND2X8TS Y A B 
.SUBCKT CLKAND2X8TS Y A B VSS VDD
X0 VDD net11 Y VDD LPPFET W=4.62U L=0.12U M=1 
X1 Y net11 VSS VSS LPNFET W=1.74U L=0.12U M=1 
X2 hnet14 B VSS VSS LPNFET W=0.74U L=0.12U M=1 
X3 net11 A hnet14 VSS LPNFET W=0.74U L=0.12U M=1 
X4 VDD B net11 VDD LPPFET W=2.06U L=0.12U M=1 
X5 VDD A net11 VDD LPPFET W=2.06U L=0.12U M=1 
.ENDS CLKAND2X8TS 

**** 
*.SUBCKT CLKBUFX12TS Y A 
.SUBCKT CLKBUFX12TS Y A VSS VDD
X0 VDD nmin Y VDD LPPFET W=7.62U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=2.82U L=0.12U M=1 
X2 VDD A nmin VDD LPPFET W=2.44U L=0.12U M=1 
X3 nmin A VSS VSS LPNFET W=0.9U L=0.12U M=1 
.ENDS CLKBUFX12TS 

**** 
*.SUBCKT CLKBUFX16TS Y A 
.SUBCKT CLKBUFX16TS Y A VSS VDD
X0 VDD nmin Y VDD LPPFET W=10.4U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=3.78U L=0.12U M=1 
X2 VDD A nmin VDD LPPFET W=3.3U L=0.12U M=1 
X3 nmin A VSS VSS LPNFET W=1.22U L=0.12U M=1 
.ENDS CLKBUFX16TS 

**** 
*.SUBCKT CLKBUFX20TS Y A 
.SUBCKT CLKBUFX20TS Y A VSS VDD
X0 VDD nmin Y VDD LPPFET W=13U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=4.74U L=0.12U M=1 
X2 VDD A nmin VDD LPPFET W=3.88U L=0.12U M=1 
X3 nmin A VSS VSS LPNFET W=1.52U L=0.12U M=1 
.ENDS CLKBUFX20TS 

**** 
*.SUBCKT CLKBUFX2TS Y A 
.SUBCKT CLKBUFX2TS Y A VSS VDD
X0 VDD nmin Y VDD LPPFET W=1.3U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=0.48U L=0.12U M=1 
X2 VDD A nmin VDD LPPFET W=0.54U L=0.12U M=1 
X3 nmin A VSS VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS CLKBUFX2TS 

**** 
*.SUBCKT CLKBUFX3TS Y A 
.SUBCKT CLKBUFX3TS Y A VSS VDD
X0 VDD nmin Y VDD LPPFET W=1.94U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=0.72U L=0.12U M=1 
X2 VDD A nmin VDD LPPFET W=0.6U L=0.12U M=1 
X3 nmin A VSS VSS LPNFET W=0.22U L=0.12U M=1 
.ENDS CLKBUFX3TS 

**** 
*.SUBCKT CLKBUFX4TS Y A 
.SUBCKT CLKBUFX4TS Y A VSS VDD
X0 VDD nmin Y VDD LPPFET W=2.54U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=0.94U L=0.12U M=1 
X2 VDD A nmin VDD LPPFET W=0.8U L=0.12U M=1 
X3 nmin A VSS VSS LPNFET W=0.3U L=0.12U M=1 
.ENDS CLKBUFX4TS 

**** 
*.SUBCKT CLKBUFX6TS Y A 
.SUBCKT CLKBUFX6TS Y A VSS VDD
X0 VDD nmin Y VDD LPPFET W=3.84U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=1.42U L=0.12U M=1 
X2 VDD A nmin VDD LPPFET W=1.16U L=0.12U M=1 
X3 nmin A VSS VSS LPNFET W=0.46U L=0.12U M=1 
.ENDS CLKBUFX6TS 

**** 
*.SUBCKT CLKBUFX8TS Y A 
.SUBCKT CLKBUFX8TS Y A VSS VDD
X0 VDD nmin Y VDD LPPFET W=5.12U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=1.84U L=0.12U M=1 
X2 VDD A nmin VDD LPPFET W=1.62U L=0.12U M=1 
X3 nmin A VSS VSS LPNFET W=0.6U L=0.12U M=1 
.ENDS CLKBUFX8TS 

**** 
*.SUBCKT CLKINVX12TS Y A 
.SUBCKT CLKINVX12TS Y A VSS VDD
X0 VDD A Y VDD LPPFET W=7.62U L=0.12U M=1 
X1 Y A VSS VSS LPNFET W=2.82U L=0.12U M=1 
.ENDS CLKINVX12TS 

**** 
*.SUBCKT CLKINVX16TS Y A 
.SUBCKT CLKINVX16TS Y A VSS VDD
X0 VDD A Y VDD LPPFET W=10.4U L=0.12U M=1 
X1 Y A VSS VSS LPNFET W=3.78U L=0.12U M=1 
.ENDS CLKINVX16TS 

**** 
*.SUBCKT CLKINVX1TS Y A 
.SUBCKT CLKINVX1TS Y A VSS VDD
X0 VDD A Y VDD LPPFET W=0.64U L=0.12U M=1 
X1 Y A VSS VSS LPNFET W=0.24U L=0.12U M=1 
.ENDS CLKINVX1TS 

**** 
*.SUBCKT CLKINVX20TS Y A 
.SUBCKT CLKINVX20TS Y A VSS VDD
X0 VDD A Y VDD LPPFET W=12.5U L=0.12U M=1 
X1 Y A VSS VSS LPNFET W=4.86U L=0.12U M=1 
.ENDS CLKINVX20TS 

**** 
*.SUBCKT CLKINVX2TS Y A 
.SUBCKT CLKINVX2TS Y A VSS VDD
X0 VDD A Y VDD LPPFET W=1.3U L=0.12U M=1 
X1 Y A VSS VSS LPNFET W=0.48U L=0.12U M=1 
.ENDS CLKINVX2TS 

**** 
*.SUBCKT CLKINVX3TS Y A 
.SUBCKT CLKINVX3TS Y A VSS VDD
X0 VDD A Y VDD LPPFET W=1.94U L=0.12U M=1 
X1 Y A VSS VSS LPNFET W=0.72U L=0.12U M=1 
.ENDS CLKINVX3TS 

**** 
*.SUBCKT CLKINVX4TS Y A 
.SUBCKT CLKINVX4TS Y A VSS VDD
X0 VDD A Y VDD LPPFET W=2.54U L=0.12U M=1 
X1 Y A VSS VSS LPNFET W=0.94U L=0.12U M=1 
.ENDS CLKINVX4TS 

**** 
*.SUBCKT CLKINVX6TS Y A 
.SUBCKT CLKINVX6TS Y A VSS VDD
X0 VDD A Y VDD LPPFET W=3.84U L=0.12U M=1 
X1 Y A VSS VSS LPNFET W=1.42U L=0.12U M=1 
.ENDS CLKINVX6TS 

**** 
*.SUBCKT CLKINVX8TS Y A 
.SUBCKT CLKINVX8TS Y A VSS VDD
X0 VDD A Y VDD LPPFET W=5.06U L=0.12U M=1 
X1 Y A VSS VSS LPNFET W=1.9U L=0.12U M=1 
.ENDS CLKINVX8TS 

**** 
*.SUBCKT CLKMX2X12TS Y A B S0 
.SUBCKT CLKMX2X12TS Y A B S0 VSS VDD
X0 net27 nmsel nmin0 VSS LPNFET W=0.38U L=0.12U M=1 
X1 net27 S0 nmin1 VSS LPNFET W=0.38U L=0.12U M=1 
X10 VDD A nmin0 VDD LPPFET W=1.02U L=0.12U M=1 
X11 nmin0 A VSS VSS LPNFET W=0.38U L=0.12U M=1 
X12 VDD B nmin1 VDD LPPFET W=1.02U L=0.12U M=1 
X13 nmin1 B VSS VSS LPNFET W=0.38U L=0.12U M=1 
X14 VDD S0 nmsel VDD LPPFET W=0.54U L=0.12U M=1 
X15 nmsel S0 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 net27 S0 nmin0 VDD LPPFET W=1.02U L=0.12U M=1 
X3 net27 nmsel nmin1 VDD LPPFET W=1.02U L=0.12U M=1 
X4 VDD net39 Y VDD LPPFET W=7.62U L=0.12U M=1 
X5 Y net39 VSS VSS LPNFET W=2.76U L=0.12U M=1 
X6 VDD net41 net39 VDD LPPFET W=3.08U L=0.12U M=1 
X7 net39 net41 VSS VSS LPNFET W=1.14U L=0.12U M=1 
X8 VDD net27 net41 VDD LPPFET W=1.24U L=0.12U M=1 
X9 net41 net27 VSS VSS LPNFET W=0.46U L=0.12U M=1 
.ENDS CLKMX2X12TS 

**** 
*.SUBCKT CLKMX2X2TS Y A B S0 
.SUBCKT CLKMX2X2TS Y A B S0 VSS VDD
X0 net25 nmsel nmin0 VSS LPNFET W=0.38U L=0.12U M=1 
X1 net25 S0 nmin1 VSS LPNFET W=0.36U L=0.12U M=1 
X10 VDD S0 nmsel VDD LPPFET W=0.54U L=0.12U M=1 
X11 nmsel S0 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 net25 S0 nmin0 VDD LPPFET W=1.02U L=0.12U M=1 
X3 net25 nmsel nmin1 VDD LPPFET W=1.02U L=0.12U M=1 
X4 VDD net25 Y VDD LPPFET W=1.28U L=0.12U M=1 
X5 Y net25 VSS VSS LPNFET W=0.48U L=0.12U M=1 
X6 VDD A nmin0 VDD LPPFET W=1.02U L=0.12U M=1 
X7 nmin0 A VSS VSS LPNFET W=0.38U L=0.12U M=1 
X8 VDD B nmin1 VDD LPPFET W=1.02U L=0.12U M=1 
X9 nmin1 B VSS VSS LPNFET W=0.36U L=0.12U M=1 
.ENDS CLKMX2X2TS 

**** 
*.SUBCKT CLKMX2X3TS Y A B S0 
.SUBCKT CLKMX2X3TS Y A B S0 VSS VDD
X0 net25 nmsel nmin0 VSS LPNFET W=0.54U L=0.12U M=1 
X1 net25 S0 nmin1 VSS LPNFET W=0.54U L=0.12U M=1 
X10 VDD S0 nmsel VDD LPPFET W=0.52U L=0.12U M=1 
X11 nmsel S0 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 net25 S0 nmin0 VDD LPPFET W=1.24U L=0.12U M=1 
X3 net25 nmsel nmin1 VDD LPPFET W=1.24U L=0.12U M=1 
X4 VDD net25 Y VDD LPPFET W=1.84U L=0.12U M=1 
X5 Y net25 VSS VSS LPNFET W=0.66U L=0.12U M=1 
X6 VDD A nmin0 VDD LPPFET W=1.24U L=0.12U M=1 
X7 nmin0 A VSS VSS LPNFET W=0.54U L=0.12U M=1 
X8 VDD B nmin1 VDD LPPFET W=1.24U L=0.12U M=1 
X9 nmin1 B VSS VSS LPNFET W=0.54U L=0.12U M=1 
.ENDS CLKMX2X3TS 

**** 
*.SUBCKT CLKMX2X4TS Y A B S0 
.SUBCKT CLKMX2X4TS Y A B S0 VSS VDD
X0 net25 nmsel nmin0 VSS LPNFET W=0.52U L=0.12U M=1 
X1 net25 S0 nmin1 VSS LPNFET W=0.44U L=0.12U M=1 
X10 VDD S0 nmsel VDD LPPFET W=0.6U L=0.12U M=1 
X11 nmsel S0 VSS VSS LPNFET W=0.22U L=0.12U M=1 
X2 net25 S0 nmin0 VDD LPPFET W=1.18U L=0.12U M=1 
X3 net25 nmsel nmin1 VDD LPPFET W=1.18U L=0.12U M=1 
X4 VDD net25 Y VDD LPPFET W=2.36U L=0.12U M=1 
X5 Y net25 VSS VSS LPNFET W=0.9U L=0.12U M=1 
X6 VDD A nmin0 VDD LPPFET W=1.18U L=0.12U M=1 
X7 nmin0 A VSS VSS LPNFET W=0.44U L=0.12U M=1 
X8 VDD B nmin1 VDD LPPFET W=1.18U L=0.12U M=1 
X9 nmin1 B VSS VSS LPNFET W=0.44U L=0.12U M=1 
.ENDS CLKMX2X4TS 

**** 
*.SUBCKT CLKMX2X6TS Y A B S0 
.SUBCKT CLKMX2X6TS Y A B S0 VSS VDD
X0 net25 nmsel nmin0 VSS LPNFET W=1.04U L=0.12U M=1 
X1 net25 S0 nmin1 VSS LPNFET W=1.04U L=0.12U M=1 
X10 VDD S0 nmsel VDD LPPFET W=1.24U L=0.12U M=1 
X11 nmsel S0 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X2 net25 S0 nmin0 VDD LPPFET W=2.82U L=0.12U M=1 
X3 net25 nmsel nmin1 VDD LPPFET W=3.06U L=0.12U M=1 
X4 VDD net25 Y VDD LPPFET W=3.84U L=0.12U M=1 
X5 Y net25 VSS VSS LPNFET W=1.42U L=0.12U M=1 
X6 VDD A nmin0 VDD LPPFET W=2.94U L=0.12U M=1 
X7 nmin0 A VSS VSS LPNFET W=1.14U L=0.12U M=1 
X8 VDD B nmin1 VDD LPPFET W=3.06U L=0.12U M=1 
X9 nmin1 B VSS VSS LPNFET W=1.12U L=0.12U M=1 
.ENDS CLKMX2X6TS 

**** 
*.SUBCKT CLKMX2X8TS Y A B S0 
.SUBCKT CLKMX2X8TS Y A B S0 VSS VDD
X0 net27 nmsel nmin0 VSS LPNFET W=0.24U L=0.12U M=1 
X1 net27 S0 nmin1 VSS LPNFET W=0.24U L=0.12U M=1 
X10 VDD A nmin0 VDD LPPFET W=0.64U L=0.12U M=1 
X11 nmin0 A VSS VSS LPNFET W=0.24U L=0.12U M=1 
X12 VDD B nmin1 VDD LPPFET W=0.64U L=0.12U M=1 
X13 nmin1 B VSS VSS LPNFET W=0.24U L=0.12U M=1 
X14 VDD S0 nmsel VDD LPPFET W=0.54U L=0.12U M=1 
X15 nmsel S0 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 net27 S0 nmin0 VDD LPPFET W=0.64U L=0.12U M=1 
X3 net27 nmsel nmin1 VDD LPPFET W=0.64U L=0.12U M=1 
X4 VDD net41 net37 VDD LPPFET W=2.06U L=0.12U M=1 
X5 net37 net41 VSS VSS LPNFET W=0.76U L=0.12U M=1 
X6 VDD net37 Y VDD LPPFET W=5.12U L=0.12U M=1 
X7 Y net37 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X8 VDD net27 net41 VDD LPPFET W=0.8U L=0.12U M=1 
X9 net41 net27 VSS VSS LPNFET W=0.3U L=0.12U M=1 
.ENDS CLKMX2X8TS 

**** 
*.SUBCKT CLKXOR2X1TS Y A B 
.SUBCKT CLKXOR2X1TS Y A B VSS VDD
X0 net29 nmin1 net37 VDD LPPFET W=0.54U L=0.12U M=1 
X1 net29 A nmin2 VDD LPPFET W=0.54U L=0.12U M=1 
X10 VDD B nmin2 VDD LPPFET W=0.6U L=0.12U M=1 
X11 nmin2 B VSS VSS LPNFET W=0.22U L=0.12U M=1 
X2 net29 A net37 VSS LPNFET W=0.2U L=0.12U M=1 
X3 net29 nmin1 nmin2 VSS LPNFET W=0.2U L=0.12U M=1 
X4 VDD net29 Y VDD LPPFET W=0.64U L=0.12U M=1 
X5 Y net29 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X6 VDD A nmin1 VDD LPPFET W=0.54U L=0.12U M=1 
X7 nmin1 A VSS VSS LPNFET W=0.2U L=0.12U M=1 
X8 VDD nmin2 net37 VDD LPPFET W=0.54U L=0.12U M=1 
X9 net37 nmin2 VSS VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS CLKXOR2X1TS 

**** 
*.SUBCKT CLKXOR2X2TS Y A B 
.SUBCKT CLKXOR2X2TS Y A B VSS VDD
X0 net29 nmin1 net37 VDD LPPFET W=0.8U L=0.12U M=1 
X1 net29 A nmin2 VDD LPPFET W=0.8U L=0.12U M=1 
X10 VDD B nmin2 VDD LPPFET W=1.08U L=0.12U M=1 
X11 nmin2 B VSS VSS LPNFET W=0.4U L=0.12U M=1 
X2 net29 A net37 VSS LPNFET W=0.3U L=0.12U M=1 
X3 net29 nmin1 nmin2 VSS LPNFET W=0.3U L=0.12U M=1 
X4 VDD net29 Y VDD LPPFET W=1.3U L=0.12U M=1 
X5 Y net29 VSS VSS LPNFET W=0.48U L=0.12U M=1 
X6 VDD A nmin1 VDD LPPFET W=0.54U L=0.12U M=1 
X7 nmin1 A VSS VSS LPNFET W=0.2U L=0.12U M=1 
X8 VDD nmin2 net37 VDD LPPFET W=0.8U L=0.12U M=1 
X9 net37 nmin2 VSS VSS LPNFET W=0.3U L=0.12U M=1 
.ENDS CLKXOR2X2TS 

**** 
*.SUBCKT CLKXOR2X4TS Y A B 
.SUBCKT CLKXOR2X4TS Y A B VSS VDD
X0 net29 nmin1 net37 VDD LPPFET W=1.5U L=0.12U M=1 
X1 net29 A nmin2 VDD LPPFET W=1.62U L=0.12U M=1 
X10 VDD B nmin2 VDD LPPFET W=2.16U L=0.12U M=1 
X11 nmin2 B VSS VSS LPNFET W=0.8U L=0.12U M=1 
X2 net29 A net37 VSS LPNFET W=0.6U L=0.12U M=1 
X3 net29 nmin1 nmin2 VSS LPNFET W=0.6U L=0.12U M=1 
X4 VDD net29 Y VDD LPPFET W=2.54U L=0.12U M=1 
X5 Y net29 VSS VSS LPNFET W=0.94U L=0.12U M=1 
X6 VDD A nmin1 VDD LPPFET W=0.54U L=0.12U M=1 
X7 nmin1 A VSS VSS LPNFET W=0.2U L=0.12U M=1 
X8 VDD nmin2 net37 VDD LPPFET W=1.5U L=0.12U M=1 
X9 net37 nmin2 VSS VSS LPNFET W=0.6U L=0.12U M=1 
.ENDS CLKXOR2X4TS 

**** 
*.SUBCKT CLKXOR2X8TS Y A B 
.SUBCKT CLKXOR2X8TS Y A B VSS VDD
X0 net29 nmin1 net37 VDD LPPFET W=3.24U L=0.12U M=1 
X1 net29 A nmin2 VDD LPPFET W=3.24U L=0.12U M=1 
X10 VDD B nmin2 VDD LPPFET W=3.88U L=0.12U M=1 
X11 nmin2 B VSS VSS LPNFET W=1.58U L=0.12U M=1 
X2 net29 A net37 VSS LPNFET W=1.2U L=0.12U M=1 
X3 net29 nmin1 nmin2 VSS LPNFET W=1.2U L=0.12U M=1 
X4 VDD net29 Y VDD LPPFET W=5.12U L=0.12U M=1 
X5 Y net29 VSS VSS LPNFET W=1.88U L=0.12U M=1 
X6 VDD A nmin1 VDD LPPFET W=1.04U L=0.12U M=1 
X7 nmin1 A VSS VSS LPNFET W=0.38U L=0.12U M=1 
X8 VDD nmin2 net37 VDD LPPFET W=3.12U L=0.12U M=1 
X9 net37 nmin2 VSS VSS LPNFET W=1.2U L=0.12U M=1 
.ENDS CLKXOR2X8TS 

**** 
*.SUBCKT CMPR22X2TS CO S A B 
.SUBCKT CMPR22X2TS CO S A B VSS VDD
X0 hnet16 A VSS VSS LPNFET W=0.48U L=0.12U M=1 
X1 net27 B hnet16 VSS LPNFET W=0.48U L=0.12U M=1 
X10 VDD B nmb VDD LPPFET W=1.02U L=0.12U M=1 
X11 nmb B VSS VSS LPNFET W=0.72U L=0.12U M=1 
X12 VDD net46 net45 VDD LPPFET W=2.56U L=0.12U M=1 
X13 net45 net46 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X14 VDD A net46 VDD LPPFET W=3.6U L=0.12U M=1 
X15 net46 A VSS VSS LPNFET W=2.58U L=0.12U M=1 
X2 VDD A net27 VDD LPPFET W=0.5U L=0.12U M=1 
X3 VDD B net27 VDD LPPFET W=0.5U L=0.12U M=1 
X4 S B net45 VDD LPPFET W=2.54U L=0.12U M=1 
X5 S nmb net46 VDD LPPFET W=2.56U L=0.12U M=1 
X6 S nmb net45 VSS LPNFET W=1.66U L=0.12U M=1 
X7 S B net46 VSS LPNFET W=1.76U L=0.12U M=1 
X8 VDD net27 CO VDD LPPFET W=1.28U L=0.12U M=1 
X9 CO net27 VSS VSS LPNFET W=0.92U L=0.12U M=1 
.ENDS CMPR22X2TS 

**** 
*.SUBCKT CMPR22X4TS CO S A B 
.SUBCKT CMPR22X4TS CO S A B VSS VDD
X0 hnet16 A VSS VSS LPNFET W=0.92U L=0.12U M=1 
X1 net27 B hnet16 VSS LPNFET W=0.92U L=0.12U M=1 
X10 VDD B nmb VDD LPPFET W=2.06U L=0.12U M=1 
X11 nmb B VSS VSS LPNFET W=1.32U L=0.12U M=1 
X12 VDD net46 net45 VDD LPPFET W=5.12U L=0.12U M=1 
X13 net45 net46 VSS VSS LPNFET W=3.68U L=0.12U M=1 
X14 VDD A net46 VDD LPPFET W=7.18U L=0.12U M=1 
X15 net46 A VSS VSS LPNFET W=4.6U L=0.12U M=1 
X2 VDD A net27 VDD LPPFET W=0.9U L=0.12U M=1 
X3 VDD B net27 VDD LPPFET W=0.9U L=0.12U M=1 
X4 S B net45 VDD LPPFET W=4.96U L=0.12U M=1 
X5 S nmb net46 VDD LPPFET W=4.96U L=0.12U M=1 
X6 S nmb net45 VSS LPNFET W=3.68U L=0.12U M=1 
X7 S B net46 VSS LPNFET W=3.68U L=0.12U M=1 
X8 VDD net27 CO VDD LPPFET W=2.56U L=0.12U M=1 
X9 CO net27 VSS VSS LPNFET W=1.84U L=0.12U M=1 
.ENDS CMPR22X4TS 

**** 
*.SUBCKT CMPR32X2TS CO S A B C 
.SUBCKT CMPR32X2TS CO S A B C VSS VDD
X0 xo nmb nma VDD LPPFET W=0.5U L=0.12U M=1 
X1 xn net109 nma VDD LPPFET W=0.5U L=0.12U M=1 
X10 xo nma net109 VSS LPNFET W=0.54U L=0.12U M=1 
X11 xn nma nmb VSS LPNFET W=0.54U L=0.12U M=1 
X12 nmcin xo net78 VSS LPNFET W=0.32U L=0.12U M=1 
X13 net78 xn nmb VSS LPNFET W=0.32U L=0.12U M=1 
X14 net108 nmcin xn VSS LPNFET W=0.34U L=0.12U M=1 
X15 net108 C xo VSS LPNFET W=0.34U L=0.12U M=1 
X16 VDD nmb net109 VDD LPPFET W=0.9U L=0.12U M=1 
X17 net109 nmb VSS VSS LPNFET W=0.64U L=0.12U M=1 
X18 VDD net108 S VDD LPPFET W=1.28U L=0.12U M=1 
X19 S net108 VSS VSS LPNFET W=0.84U L=0.12U M=1 
X2 xn nma net109 VDD LPPFET W=0.76U L=0.12U M=1 
X20 VDD net78 CO VDD LPPFET W=1.28U L=0.12U M=1 
X21 CO net78 VSS VSS LPNFET W=0.84U L=0.12U M=1 
X22 VDD C nmcin VDD LPPFET W=0.5U L=0.12U M=1 
X23 nmcin C VSS VSS LPNFET W=0.32U L=0.12U M=1 
X24 VDD B nmb VDD LPPFET W=1.28U L=0.12U M=1 
X25 nmb B VSS VSS LPNFET W=0.92U L=0.12U M=1 
X26 VDD A nma VDD LPPFET W=1.28U L=0.12U M=1 
X27 nma A VSS VSS LPNFET W=0.92U L=0.12U M=1 
X3 xo nma nmb VDD LPPFET W=0.76U L=0.12U M=1 
X4 nmcin xn net78 VDD LPPFET W=0.5U L=0.12U M=1 
X5 net78 xo nmb VDD LPPFET W=0.5U L=0.12U M=1 
X6 net108 C xn VDD LPPFET W=0.5U L=0.12U M=1 
X7 net108 nmcin xo VDD LPPFET W=0.5U L=0.12U M=1 
X8 xo net109 nma VSS LPNFET W=0.34U L=0.12U M=1 
X9 xn nmb nma VSS LPNFET W=0.34U L=0.12U M=1 
.ENDS CMPR32X2TS 

**** 
*.SUBCKT CMPR32X4TS CO S A B C 
.SUBCKT CMPR32X4TS CO S A B C VSS VDD
X0 xo nmb nma VDD LPPFET W=0.5U L=0.12U M=1 
X1 xn net111 nma VDD LPPFET W=0.5U L=0.12U M=1 
X10 xo nma net111 VSS LPNFET W=0.54U L=0.12U M=1 
X11 xn nma nmb VSS LPNFET W=0.54U L=0.12U M=1 
X12 nmcin xo net80 VSS LPNFET W=0.32U L=0.12U M=1 
X13 net80 xn nmb VSS LPNFET W=0.32U L=0.12U M=1 
X14 net110 nmcin xn VSS LPNFET W=0.36U L=0.12U M=1 
X15 net110 C xo VSS LPNFET W=0.36U L=0.12U M=1 
X16 VDD nmb net111 VDD LPPFET W=0.9U L=0.12U M=1 
X17 net111 nmb VSS VSS LPNFET W=0.64U L=0.12U M=1 
X18 VDD net110 S VDD LPPFET W=2.56U L=0.12U M=1 
X19 S net110 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X2 xn nma net111 VDD LPPFET W=0.76U L=0.12U M=1 
X20 VDD net80 CO VDD LPPFET W=2.56U L=0.12U M=1 
X21 CO net80 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X22 VDD C nmcin VDD LPPFET W=0.5U L=0.12U M=1 
X23 nmcin C VSS VSS LPNFET W=0.36U L=0.12U M=1 
X24 VDD B nmb VDD LPPFET W=1.28U L=0.12U M=1 
X25 nmb B VSS VSS LPNFET W=0.92U L=0.12U M=1 
X26 VDD A nma VDD LPPFET W=1.28U L=0.12U M=1 
X27 nma A VSS VSS LPNFET W=0.92U L=0.12U M=1 
X3 xo nma nmb VDD LPPFET W=0.76U L=0.12U M=1 
X4 nmcin xn net80 VDD LPPFET W=0.5U L=0.12U M=1 
X5 net80 xo nmb VDD LPPFET W=0.5U L=0.12U M=1 
X6 net110 C xn VDD LPPFET W=0.5U L=0.12U M=1 
X7 net110 nmcin xo VDD LPPFET W=0.5U L=0.12U M=1 
X8 xo net111 nma VSS LPNFET W=0.34U L=0.12U M=1 
X9 xn nmb nma VSS LPNFET W=0.34U L=0.12U M=1 
.ENDS CMPR32X4TS 

**** 
*.SUBCKT CMPR42X1TS CO ICO S A B C D ICI 
.SUBCKT CMPR42X1TS CO ICO S A B C D ICI VSS VDD
X0 net92 net90 nmin3 VSS LPNFET W=0.36U L=0.12U M=1 
X1 net92 net144 nmcin VSS LPNFET W=0.36U L=0.12U M=1 
X10 net125 D nmin2 VSS LPNFET W=0.56U L=0.12U M=1 
X11 net125 nmin3 net128 VSS LPNFET W=0.56U L=0.12U M=1 
X12 net128 nmin2 VSS VSS LPNFET W=0.56U L=0.12U M=1 
X13 net144 net133 net125 VSS LPNFET W=0.56U L=0.12U M=1 
X14 net144 net125 net133 VSS LPNFET W=0.56U L=0.12U M=1 
X15 net140 net90 nmcin VSS LPNFET W=0.36U L=0.12U M=1 
X16 net140 net144 net143 VSS LPNFET W=0.36U L=0.12U M=1 
X17 net143 nmcin VSS VSS LPNFET W=0.36U L=0.12U M=1 
X18 net92 net144 nmin3 VDD LPPFET W=0.5U L=0.12U M=1 
X19 net92 net90 nmcin VDD LPPFET W=0.5U L=0.12U M=1 
X2 nmco B net101 VSS LPNFET W=0.36U L=0.12U M=1 
X20 net154 A VDD VDD LPPFET W=0.5U L=0.12U M=1 
X21 nmco B net154 VDD LPPFET W=0.5U L=0.12U M=1 
X22 nmco C net161 VDD LPPFET W=0.5U L=0.12U M=1 
X23 net161 B VDD VDD LPPFET W=0.5U L=0.12U M=1 
X24 net161 A VDD VDD LPPFET W=0.5U L=0.12U M=1 
X25 net183 nmin1 nmin0 VDD LPPFET W=0.78U L=0.12U M=1 
X26 net183 B net173 VDD LPPFET W=0.78U L=0.12U M=1 
X27 net173 nmin0 VDD VDD LPPFET W=0.78U L=0.12U M=1 
X28 net125 nmin3 nmin2 VDD LPPFET W=0.78U L=0.12U M=1 
X29 net125 D net182 VDD LPPFET W=0.78U L=0.12U M=1 
X3 net101 A VSS VSS LPNFET W=0.36U L=0.12U M=1 
X30 net182 nmin2 VDD VDD LPPFET W=0.78U L=0.12U M=1 
X31 net144 net183 net125 VDD LPPFET W=0.78U L=0.12U M=1 
X32 net144 net125 net183 VDD LPPFET W=0.78U L=0.12U M=1 
X33 net140 net144 nmcin VDD LPPFET W=0.5U L=0.12U M=1 
X34 net140 net90 net193 VDD LPPFET W=0.5U L=0.12U M=1 
X35 net193 nmcin VDD VDD LPPFET W=0.5U L=0.12U M=1 
X36 VDD nmco ICO VDD LPPFET W=0.64U L=0.12U M=1 
X37 ICO nmco VSS VSS LPNFET W=0.46U L=0.12U M=1 
X38 VDD net92 CO VDD LPPFET W=0.64U L=0.12U M=1 
X39 CO net92 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X4 net104 B VSS VSS LPNFET W=0.36U L=0.12U M=1 
X40 VDD net183 net133 VDD LPPFET W=0.78U L=0.12U M=1 
X41 net133 net183 VSS VSS LPNFET W=0.54U L=0.12U M=1 
X42 VDD A nmin0 VDD LPPFET W=0.78U L=0.12U M=1 
X43 nmin0 A VSS VSS LPNFET W=0.56U L=0.12U M=1 
X44 VDD B nmin1 VDD LPPFET W=0.28U L=0.12U M=1 
X45 nmin1 B VSS VSS LPNFET W=0.2U L=0.12U M=1 
X46 VDD C nmin2 VDD LPPFET W=0.78U L=0.12U M=1 
X47 nmin2 C VSS VSS LPNFET W=0.56U L=0.12U M=1 
X48 VDD D nmin3 VDD LPPFET W=0.84U L=0.12U M=1 
X49 nmin3 D VSS VSS LPNFET W=0.6U L=0.12U M=1 
X5 net104 A VSS VSS LPNFET W=0.36U L=0.12U M=1 
X50 VDD net144 net90 VDD LPPFET W=0.3U L=0.12U M=1 
X51 net90 net144 VSS VSS LPNFET W=0.22U L=0.12U M=1 
X52 VDD ICI nmcin VDD LPPFET W=0.68U L=0.12U M=1 
X53 nmcin ICI VSS VSS LPNFET W=0.52U L=0.12U M=1 
X54 VDD net140 S VDD LPPFET W=0.64U L=0.12U M=1 
X55 S net140 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X6 nmco C net104 VSS LPNFET W=0.36U L=0.12U M=1 
X7 net183 B nmin0 VSS LPNFET W=0.56U L=0.12U M=1 
X8 net183 nmin1 net119 VSS LPNFET W=0.56U L=0.12U M=1 
X9 net119 nmin0 VSS VSS LPNFET W=0.56U L=0.12U M=1 
.ENDS CMPR42X1TS 

**** 
*.SUBCKT CMPR42X2TS CO ICO S A B C D ICI 
.SUBCKT CMPR42X2TS CO ICO S A B C D ICI VSS VDD
X0 net92 net90 nmin3 VSS LPNFET W=0.74U L=0.12U M=1 
X1 net92 net144 nmcin VSS LPNFET W=0.74U L=0.12U M=1 
X10 net125 D nmin2 VSS LPNFET W=0.84U L=0.12U M=1 
X11 net125 nmin3 net128 VSS LPNFET W=0.84U L=0.12U M=1 
X12 net128 nmin2 VSS VSS LPNFET W=0.84U L=0.12U M=1 
X13 net144 net133 net125 VSS LPNFET W=0.9U L=0.12U M=1 
X14 net144 net125 net133 VSS LPNFET W=0.9U L=0.12U M=1 
X15 net140 net90 nmcin VSS LPNFET W=0.74U L=0.12U M=1 
X16 net140 net144 net143 VSS LPNFET W=0.74U L=0.12U M=1 
X17 net143 nmcin VSS VSS LPNFET W=0.74U L=0.12U M=1 
X18 net92 net144 nmin3 VDD LPPFET W=1.02U L=0.12U M=1 
X19 net92 net90 nmcin VDD LPPFET W=1.02U L=0.12U M=1 
X2 nmco B net97 VSS LPNFET W=0.74U L=0.12U M=1 
X20 net154 A VDD VDD LPPFET W=1.02U L=0.12U M=1 
X21 nmco B net154 VDD LPPFET W=1.02U L=0.12U M=1 
X22 nmco C net161 VDD LPPFET W=1.02U L=0.12U M=1 
X23 net161 B VDD VDD LPPFET W=1.02U L=0.12U M=1 
X24 net161 A VDD VDD LPPFET W=1.02U L=0.12U M=1 
X25 net183 nmin1 nmin0 VDD LPPFET W=1.16U L=0.12U M=1 
X26 net183 B net169 VDD LPPFET W=1.16U L=0.12U M=1 
X27 net169 nmin0 VDD VDD LPPFET W=1.16U L=0.12U M=1 
X28 net125 nmin3 nmin2 VDD LPPFET W=1.16U L=0.12U M=1 
X29 net125 D net178 VDD LPPFET W=1.26U L=0.12U M=1 
X3 net97 A VSS VSS LPNFET W=0.74U L=0.12U M=1 
X30 net178 nmin2 VDD VDD LPPFET W=1.26U L=0.12U M=1 
X31 net144 net183 net125 VDD LPPFET W=1.16U L=0.12U M=1 
X32 net144 net125 net183 VDD LPPFET W=1.16U L=0.12U M=1 
X33 net140 net144 nmcin VDD LPPFET W=1U L=0.12U M=1 
X34 net140 net90 net197 VDD LPPFET W=1U L=0.12U M=1 
X35 net197 nmcin VDD VDD LPPFET W=1U L=0.12U M=1 
X36 VDD nmco ICO VDD LPPFET W=1.28U L=0.12U M=1 
X37 ICO nmco VSS VSS LPNFET W=0.92U L=0.12U M=1 
X38 VDD net92 CO VDD LPPFET W=1.28U L=0.12U M=1 
X39 CO net92 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X4 net104 B VSS VSS LPNFET W=0.74U L=0.12U M=1 
X40 VDD net183 net133 VDD LPPFET W=1.16U L=0.12U M=1 
X41 net133 net183 VSS VSS LPNFET W=0.9U L=0.12U M=1 
X42 VDD A nmin0 VDD LPPFET W=1.16U L=0.12U M=1 
X43 nmin0 A VSS VSS LPNFET W=0.72U L=0.12U M=1 
X44 VDD B nmin1 VDD LPPFET W=0.38U L=0.12U M=1 
X45 nmin1 B VSS VSS LPNFET W=0.28U L=0.12U M=1 
X46 VDD C nmin2 VDD LPPFET W=1.16U L=0.12U M=1 
X47 nmin2 C VSS VSS LPNFET W=0.92U L=0.12U M=1 
X48 VDD D nmin3 VDD LPPFET W=1.16U L=0.12U M=1 
X49 nmin3 D VSS VSS LPNFET W=0.92U L=0.12U M=1 
X5 net104 A VSS VSS LPNFET W=0.74U L=0.12U M=1 
X50 VDD net144 net90 VDD LPPFET W=0.64U L=0.12U M=1 
X51 net90 net144 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X52 VDD ICI nmcin VDD LPPFET W=1.28U L=0.12U M=1 
X53 nmcin ICI VSS VSS LPNFET W=0.82U L=0.12U M=1 
X54 VDD net140 S VDD LPPFET W=1.26U L=0.12U M=1 
X55 S net140 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X6 nmco C net104 VSS LPNFET W=0.74U L=0.12U M=1 
X7 net183 B nmin0 VSS LPNFET W=0.92U L=0.12U M=1 
X8 net183 nmin1 net119 VSS LPNFET W=0.9U L=0.12U M=1 
X9 net119 nmin0 VSS VSS LPNFET W=0.9U L=0.12U M=1 
.ENDS CMPR42X2TS 

**** 
*.SUBCKT CMPR42X4TS CO ICO S A B C D ICI 
.SUBCKT CMPR42X4TS CO ICO S A B C D ICI VSS VDD
X0 net99 nmcin VSS VSS LPNFET W=0.74U L=0.12U M=1 
X1 net100 net173 net99 VSS LPNFET W=0.74U L=0.12U M=1 
X10 nmco C net121 VSS LPNFET W=1.34U L=0.12U M=1 
X11 net212 B nmin0 VSS LPNFET W=0.92U L=0.12U M=1 
X12 net212 nmin1 net132 VSS LPNFET W=0.86U L=0.12U M=1 
X13 net132 nmin0 VSS VSS LPNFET W=0.86U L=0.12U M=1 
X14 net142 D nmin2 VSS LPNFET W=0.86U L=0.12U M=1 
X15 net142 nmin3 net145 VSS LPNFET W=0.92U L=0.12U M=1 
X16 net145 nmin2 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X17 net173 net150 net142 VSS LPNFET W=0.86U L=0.12U M=1 
X18 net173 net142 net150 VSS LPNFET W=0.86U L=0.12U M=1 
X19 net100 net107 nmcin VSS LPNFET W=1.54U L=0.12U M=1 
X2 net105 A VSS VSS LPNFET W=0.74U L=0.12U M=1 
X20 net100 net173 net160 VSS LPNFET W=0.74U L=0.12U M=1 
X21 net160 nmcin VSS VSS LPNFET W=0.74U L=0.12U M=1 
X22 net100 net107 net166 VDD LPPFET W=0.8U L=0.12U M=1 
X23 net166 nmcin VDD VDD LPPFET W=0.8U L=0.12U M=1 
X24 nmco B net172 VDD LPPFET W=1.02U L=0.12U M=1 
X25 net172 A VDD VDD LPPFET W=1.02U L=0.12U M=1 
X26 net109 net173 nmin3 VDD LPPFET W=2.06U L=0.12U M=1 
X27 net109 net107 nmcin VDD LPPFET W=2.04U L=0.12U M=1 
X28 net183 A VDD VDD LPPFET W=1.02U L=0.12U M=1 
X29 nmco B net183 VDD LPPFET W=1.02U L=0.12U M=1 
X3 nmco B net105 VSS LPNFET W=0.74U L=0.12U M=1 
X30 nmco C net190 VDD LPPFET W=1.92U L=0.12U M=1 
X31 net190 B VDD VDD LPPFET W=2.04U L=0.12U M=1 
X32 net190 A VDD VDD LPPFET W=2.04U L=0.12U M=1 
X33 net212 nmin1 nmin0 VDD LPPFET W=1.16U L=0.12U M=1 
X34 net212 B net202 VDD LPPFET W=1.16U L=0.12U M=1 
X35 net202 nmin0 VDD VDD LPPFET W=1.16U L=0.12U M=1 
X36 net142 nmin3 nmin2 VDD LPPFET W=1.16U L=0.12U M=1 
X37 net142 D net211 VDD LPPFET W=1.16U L=0.12U M=1 
X38 net211 nmin2 VDD VDD LPPFET W=1.16U L=0.12U M=1 
X39 net173 net212 net142 VDD LPPFET W=1.16U L=0.12U M=1 
X4 net109 net107 nmin3 VSS LPNFET W=1.34U L=0.12U M=1 
X40 net173 net142 net212 VDD LPPFET W=1.16U L=0.12U M=1 
X41 net100 net173 nmcin VDD LPPFET W=1.92U L=0.12U M=1 
X42 net100 net107 net222 VDD LPPFET W=0.8U L=0.12U M=1 
X43 net222 nmcin VDD VDD LPPFET W=0.8U L=0.12U M=1 
X44 VDD nmco ICO VDD LPPFET W=2.56U L=0.12U M=1 
X45 ICO nmco VSS VSS LPNFET W=1.8U L=0.12U M=1 
X46 VDD net109 CO VDD LPPFET W=2.56U L=0.12U M=1 
X47 CO net109 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X48 VDD net212 net150 VDD LPPFET W=1.16U L=0.12U M=1 
X49 net150 net212 VSS VSS LPNFET W=0.86U L=0.12U M=1 
X5 net109 net173 nmcin VSS LPNFET W=1.48U L=0.12U M=1 
X50 VDD A nmin0 VDD LPPFET W=1.16U L=0.12U M=1 
X51 nmin0 A VSS VSS LPNFET W=0.72U L=0.12U M=1 
X52 VDD B nmin1 VDD LPPFET W=0.38U L=0.12U M=1 
X53 nmin1 B VSS VSS LPNFET W=0.3U L=0.12U M=1 
X54 VDD C nmin2 VDD LPPFET W=1.16U L=0.12U M=1 
X55 nmin2 C VSS VSS LPNFET W=0.86U L=0.12U M=1 
X56 VDD D nmin3 VDD LPPFET W=1.16U L=0.12U M=1 
X57 nmin3 D VSS VSS LPNFET W=0.86U L=0.12U M=1 
X58 VDD net173 net107 VDD LPPFET W=1.24U L=0.12U M=1 
X59 net107 net173 VSS VSS LPNFET W=0.9U L=0.12U M=1 
X6 nmco B net118 VSS LPNFET W=0.74U L=0.12U M=1 
X60 VDD ICI nmcin VDD LPPFET W=1.24U L=0.12U M=1 
X61 nmcin ICI VSS VSS LPNFET W=0.9U L=0.12U M=1 
X62 VDD net100 S VDD LPPFET W=2.56U L=0.12U M=1 
X63 S net100 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X7 net118 A VSS VSS LPNFET W=0.74U L=0.12U M=1 
X8 net121 B VSS VSS LPNFET W=1.44U L=0.12U M=1 
X9 net121 A VSS VSS LPNFET W=1.48U L=0.12U M=1 
.ENDS CMPR42X4TS 

**** 
*.SUBCKT DFFHQX1TS Q CK D 
.SUBCKT DFFHQX1TS Q CK D VSS VDD
X0 VDD c hnet20 VDD LPPFET W=0.58U L=0.12U M=1 
X1 hnet20 nmin pm VDD LPPFET W=0.58U L=0.12U M=1 
X10 pm c hnet26 VSS LPNFET W=0.2U L=0.12U M=1 
X11 hnet28 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X12 VDD m hnet28 VDD LPPFET W=0.28U L=0.12U M=1 
X13 hnet32 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X14 net73 cn hnet32 VSS LPNFET W=0.2U L=0.12U M=1 
X15 hnet34 c net73 VDD LPPFET W=0.26U L=0.12U M=1 
X16 VDD s hnet34 VDD LPPFET W=0.26U L=0.12U M=1 
X17 VDD D nmin VDD LPPFET W=0.28U L=0.12U M=1 
X18 nmin D VSS VSS LPNFET W=0.2U L=0.12U M=1 
X19 VDD pm m VDD LPPFET W=0.96U L=0.12U M=1 
X2 hnet24 cn VSS VSS LPNFET W=0.42U L=0.12U M=1 
X20 m pm VSS VSS LPNFET W=0.5U L=0.12U M=1 
X21 VDD net73 s VDD LPPFET W=0.28U L=0.12U M=1 
X22 s net73 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X23 VDD net73 Q VDD LPPFET W=0.74U L=0.12U M=1 
X24 Q net73 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X25 VDD net86 c VDD LPPFET W=0.84U L=0.12U M=1 
X26 c net86 VSS VSS LPNFET W=0.3U L=0.12U M=1 
X27 VDD CK net86 VDD LPPFET W=0.28U L=0.12U M=1 
X28 net86 CK VSS VSS LPNFET W=0.28U L=0.12U M=1 
X3 pm nmin hnet24 VSS LPNFET W=0.42U L=0.12U M=1 
X4 net57 CK VDD VDD LPPFET W=0.7U L=0.12U M=1 
X5 cn c net57 VDD LPPFET W=0.5U L=0.12U M=1 
X6 net73 cn m VDD LPPFET W=0.96U L=0.12U M=1 
X7 cn CK VSS VSS LPNFET W=0.2U L=0.12U M=1 
X8 net73 c m VSS LPNFET W=0.48U L=0.12U M=1 
X9 hnet26 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS DFFHQX1TS 

**** 
*.SUBCKT DFFHQX2TS Q CK D 
.SUBCKT DFFHQX2TS Q CK D VSS VDD
X0 VDD c hnet20 VDD LPPFET W=1U L=0.12U M=1 
X1 hnet20 nmin pm VDD LPPFET W=1U L=0.12U M=1 
X10 pm c hnet26 VSS LPNFET W=0.2U L=0.12U M=1 
X11 hnet28 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X12 VDD m hnet28 VDD LPPFET W=0.28U L=0.12U M=1 
X13 hnet32 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X14 net73 cn hnet32 VSS LPNFET W=0.2U L=0.12U M=1 
X15 hnet34 c net73 VDD LPPFET W=0.28U L=0.12U M=1 
X16 VDD s hnet34 VDD LPPFET W=0.28U L=0.12U M=1 
X17 VDD D nmin VDD LPPFET W=0.34U L=0.12U M=1 
X18 nmin D VSS VSS LPNFET W=0.24U L=0.12U M=1 
X19 VDD pm m VDD LPPFET W=1.56U L=0.12U M=1 
X2 hnet24 cn VSS VSS LPNFET W=0.68U L=0.12U M=1 
X20 m pm VSS VSS LPNFET W=0.86U L=0.12U M=1 
X21 VDD net73 s VDD LPPFET W=0.28U L=0.12U M=1 
X22 s net73 VSS VSS LPNFET W=0.18U L=0.12U M=1 
X23 VDD net73 Q VDD LPPFET W=1.3U L=0.12U M=1 
X24 Q net73 VSS VSS LPNFET W=0.88U L=0.12U M=1 
X25 VDD net86 c VDD LPPFET W=1.18U L=0.12U M=1 
X26 c net86 VSS VSS LPNFET W=0.42U L=0.12U M=1 
X27 VDD CK net86 VDD LPPFET W=0.32U L=0.12U M=1 
X28 net86 CK VSS VSS LPNFET W=0.32U L=0.12U M=1 
X3 pm nmin hnet24 VSS LPNFET W=0.68U L=0.12U M=1 
X4 net55 CK VDD VDD LPPFET W=0.9U L=0.12U M=1 
X5 cn c net55 VDD LPPFET W=0.68U L=0.12U M=1 
X6 net73 cn m VDD LPPFET W=1.56U L=0.12U M=1 
X7 cn CK VSS VSS LPNFET W=0.26U L=0.12U M=1 
X8 net73 c m VSS LPNFET W=0.82U L=0.12U M=1 
X9 hnet26 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS DFFHQX2TS 

**** 
*.SUBCKT DFFHQX4TS Q CK D 
.SUBCKT DFFHQX4TS Q CK D VSS VDD
X0 hnet21 cn VSS VSS LPNFET W=0.6U L=0.12U M=1 
X1 pm nmin hnet21 VSS LPNFET W=0.6U L=0.12U M=1 
X10 net73 cn m VDD LPPFET W=2.82U L=0.12U M=1 
X11 cn CK VSS VSS LPNFET W=0.48U L=0.12U M=1 
X12 net73 c m VSS LPNFET W=1.4U L=0.12U M=1 
X13 hnet28 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X14 pm c hnet28 VSS LPNFET W=0.2U L=0.12U M=1 
X15 hnet30 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X16 VDD m hnet30 VDD LPPFET W=0.28U L=0.12U M=1 
X17 hnet34 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X18 net73 cn hnet34 VSS LPNFET W=0.2U L=0.12U M=1 
X19 hnet36 c net73 VDD LPPFET W=0.28U L=0.12U M=1 
X2 hnet17 cn VSS VSS LPNFET W=0.6U L=0.12U M=1 
X20 VDD s hnet36 VDD LPPFET W=0.28U L=0.12U M=1 
X21 VDD D nmin VDD LPPFET W=0.62U L=0.12U M=1 
X22 nmin D VSS VSS LPNFET W=0.44U L=0.12U M=1 
X23 VDD pm m VDD LPPFET W=2.56U L=0.12U M=1 
X24 m pm VSS VSS LPNFET W=1.56U L=0.12U M=1 
X25 VDD net73 s VDD LPPFET W=0.28U L=0.12U M=1 
X26 s net73 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X27 VDD net73 Q VDD LPPFET W=2.6U L=0.12U M=1 
X28 Q net73 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X29 VDD net86 c VDD LPPFET W=1.92U L=0.12U M=1 
X3 pm nmin hnet17 VSS LPNFET W=0.6U L=0.12U M=1 
X30 c net86 VSS VSS LPNFET W=0.72U L=0.12U M=1 
X31 VDD CK net86 VDD LPPFET W=0.54U L=0.12U M=1 
X32 net86 CK VSS VSS LPNFET W=0.54U L=0.12U M=1 
X4 VDD c hnet26 VDD LPPFET W=0.88U L=0.12U M=1 
X5 hnet26 nmin pm VDD LPPFET W=0.88U L=0.12U M=1 
X6 VDD c hnet23 VDD LPPFET W=0.88U L=0.12U M=1 
X7 hnet23 nmin pm VDD LPPFET W=0.88U L=0.12U M=1 
X8 net57 CK VDD VDD LPPFET W=1.3U L=0.12U M=1 
X9 cn c net57 VDD LPPFET W=1.3U L=0.12U M=1 
.ENDS DFFHQX4TS 

**** 
*.SUBCKT DFFHQX8TS Q CK D 
.SUBCKT DFFHQX8TS Q CK D VSS VDD
X0 hnet21 cn VSS VSS LPNFET W=0.6U L=0.12U M=1 
X1 pm nmin hnet21 VSS LPNFET W=0.6U L=0.12U M=1 
X10 net73 cn m VDD LPPFET W=2.82U L=0.12U M=1 
X11 cn CK VSS VSS LPNFET W=0.48U L=0.12U M=1 
X12 net73 c m VSS LPNFET W=1.4U L=0.12U M=1 
X13 hnet28 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X14 pm c hnet28 VSS LPNFET W=0.2U L=0.12U M=1 
X15 hnet30 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X16 VDD m hnet30 VDD LPPFET W=0.28U L=0.12U M=1 
X17 hnet34 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X18 net73 cn hnet34 VSS LPNFET W=0.2U L=0.12U M=1 
X19 hnet36 c net73 VDD LPPFET W=0.28U L=0.12U M=1 
X2 hnet17 cn VSS VSS LPNFET W=0.6U L=0.12U M=1 
X20 VDD s hnet36 VDD LPPFET W=0.28U L=0.12U M=1 
X21 VDD D nmin VDD LPPFET W=0.62U L=0.12U M=1 
X22 nmin D VSS VSS LPNFET W=0.44U L=0.12U M=1 
X23 VDD pm m VDD LPPFET W=2.56U L=0.12U M=1 
X24 m pm VSS VSS LPNFET W=1.56U L=0.12U M=1 
X25 VDD net73 s VDD LPPFET W=0.28U L=0.12U M=1 
X26 s net73 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X27 VDD net73 Q VDD LPPFET W=5.9U L=0.12U M=1 
X28 Q net73 VSS VSS LPNFET W=3.7U L=0.12U M=1 
X29 VDD net86 c VDD LPPFET W=1.92U L=0.12U M=1 
X3 pm nmin hnet17 VSS LPNFET W=0.6U L=0.12U M=1 
X30 c net86 VSS VSS LPNFET W=0.72U L=0.12U M=1 
X31 VDD CK net86 VDD LPPFET W=0.54U L=0.12U M=1 
X32 net86 CK VSS VSS LPNFET W=0.54U L=0.12U M=1 
X4 VDD c hnet26 VDD LPPFET W=0.88U L=0.12U M=1 
X5 hnet26 nmin pm VDD LPPFET W=0.88U L=0.12U M=1 
X6 VDD c hnet23 VDD LPPFET W=0.88U L=0.12U M=1 
X7 hnet23 nmin pm VDD LPPFET W=0.88U L=0.12U M=1 
X8 net57 CK VDD VDD LPPFET W=1.3U L=0.12U M=1 
X9 cn c net57 VDD LPPFET W=1.3U L=0.12U M=1 
.ENDS DFFHQX8TS 

**** 
*.SUBCKT DFFNSRX1TS Q QN CKN D RN SN 
.SUBCKT DFFNSRX1TS Q QN CKN D RN SN VSS VDD
X0 m SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X1 m pm net63 VDD LPPFET W=0.42U L=0.12U M=1 
X10 net96 s net94 VSS LPNFET W=0.2U L=0.12U M=1 
X11 net94 SN VSS VSS LPNFET W=0.4U L=0.12U M=1 
X12 net100 cn net96 VSS LPNFET W=0.2U L=0.12U M=1 
X13 net100 c m VSS LPNFET W=0.2U L=0.12U M=1 
X14 hnet24 D VSS VSS LPNFET W=0.2U L=0.12U M=1 
X15 pm cn hnet24 VSS LPNFET W=0.2U L=0.12U M=1 
X16 hnet26 c pm VDD LPPFET W=0.28U L=0.12U M=1 
X17 VDD D hnet26 VDD LPPFET W=0.28U L=0.12U M=1 
X18 hnet30 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X19 pm c hnet30 VSS LPNFET W=0.2U L=0.12U M=1 
X2 net63 net113 VDD VDD LPPFET W=0.56U L=0.12U M=1 
X20 hnet32 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X21 VDD m hnet32 VDD LPPFET W=0.28U L=0.12U M=1 
X22 VDD s net109 VDD LPPFET W=0.28U L=0.12U M=1 
X23 net109 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X24 VDD s Q VDD LPPFET W=0.64U L=0.12U M=1 
X25 Q s VSS VSS LPNFET W=0.46U L=0.12U M=1 
X26 VDD RN net113 VDD LPPFET W=0.28U L=0.12U M=1 
X27 net113 RN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X28 VDD net100 s VDD LPPFET W=0.28U L=0.12U M=1 
X29 s net100 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 net100 SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X30 VDD net109 QN VDD LPPFET W=0.64U L=0.12U M=1 
X31 QN net109 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X32 VDD CKN c VDD LPPFET W=0.42U L=0.12U M=1 
X33 c CKN VSS VSS LPNFET W=0.3U L=0.12U M=1 
X34 VDD c cn VDD LPPFET W=0.28U L=0.12U M=1 
X35 cn c VSS VSS LPNFET W=0.2U L=0.12U M=1 
X4 net73 s net63 VDD LPPFET W=0.28U L=0.12U M=1 
X5 net100 c net73 VDD LPPFET W=0.28U L=0.12U M=1 
X6 net100 cn m VDD LPPFET W=0.28U L=0.12U M=1 
X7 m net113 net94 VSS LPNFET W=0.2U L=0.12U M=1 
X8 m pm net94 VSS LPNFET W=0.3U L=0.12U M=1 
X9 net100 net113 net94 VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS DFFNSRX1TS 

**** 
*.SUBCKT DFFNSRX2TS Q QN CKN D RN SN 
.SUBCKT DFFNSRX2TS Q QN CKN D RN SN VSS VDD
X0 m SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X1 m pm net63 VDD LPPFET W=0.42U L=0.12U M=1 
X10 net96 s net94 VSS LPNFET W=0.2U L=0.12U M=1 
X11 net94 SN VSS VSS LPNFET W=0.4U L=0.12U M=1 
X12 net100 cn net96 VSS LPNFET W=0.2U L=0.12U M=1 
X13 net100 c m VSS LPNFET W=0.2U L=0.12U M=1 
X14 hnet24 D VSS VSS LPNFET W=0.2U L=0.12U M=1 
X15 pm cn hnet24 VSS LPNFET W=0.2U L=0.12U M=1 
X16 hnet26 c pm VDD LPPFET W=0.28U L=0.12U M=1 
X17 VDD D hnet26 VDD LPPFET W=0.28U L=0.12U M=1 
X18 hnet30 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X19 pm c hnet30 VSS LPNFET W=0.2U L=0.12U M=1 
X2 net63 net113 VDD VDD LPPFET W=0.56U L=0.12U M=1 
X20 hnet32 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X21 VDD m hnet32 VDD LPPFET W=0.28U L=0.12U M=1 
X22 VDD s net109 VDD LPPFET W=0.3U L=0.12U M=1 
X23 net109 s VSS VSS LPNFET W=0.22U L=0.12U M=1 
X24 VDD s Q VDD LPPFET W=1.28U L=0.12U M=1 
X25 Q s VSS VSS LPNFET W=0.92U L=0.12U M=1 
X26 VDD RN net113 VDD LPPFET W=0.28U L=0.12U M=1 
X27 net113 RN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X28 VDD net100 s VDD LPPFET W=0.34U L=0.12U M=1 
X29 s net100 VSS VSS LPNFET W=0.26U L=0.12U M=1 
X3 net100 SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X30 VDD net109 QN VDD LPPFET W=1.28U L=0.12U M=1 
X31 QN net109 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X32 VDD CKN c VDD LPPFET W=0.42U L=0.12U M=1 
X33 c CKN VSS VSS LPNFET W=0.3U L=0.12U M=1 
X34 VDD c cn VDD LPPFET W=0.28U L=0.12U M=1 
X35 cn c VSS VSS LPNFET W=0.2U L=0.12U M=1 
X4 net73 s net63 VDD LPPFET W=0.28U L=0.12U M=1 
X5 net100 c net73 VDD LPPFET W=0.28U L=0.12U M=1 
X6 net100 cn m VDD LPPFET W=0.28U L=0.12U M=1 
X7 m net113 net94 VSS LPNFET W=0.2U L=0.12U M=1 
X8 m pm net94 VSS LPNFET W=0.3U L=0.12U M=1 
X9 net100 net113 net94 VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS DFFNSRX2TS 

**** 
*.SUBCKT DFFNSRX4TS Q QN CKN D RN SN 
.SUBCKT DFFNSRX4TS Q QN CKN D RN SN VSS VDD
X0 m SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X1 m pm net63 VDD LPPFET W=0.46U L=0.12U M=1 
X10 net96 s net94 VSS LPNFET W=0.2U L=0.12U M=1 
X11 net94 SN VSS VSS LPNFET W=0.46U L=0.12U M=1 
X12 net100 cn net96 VSS LPNFET W=0.2U L=0.12U M=1 
X13 net100 c m VSS LPNFET W=0.22U L=0.12U M=1 
X14 hnet24 D VSS VSS LPNFET W=0.2U L=0.12U M=1 
X15 pm cn hnet24 VSS LPNFET W=0.2U L=0.12U M=1 
X16 hnet26 c pm VDD LPPFET W=0.28U L=0.12U M=1 
X17 VDD D hnet26 VDD LPPFET W=0.28U L=0.12U M=1 
X18 hnet30 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X19 pm c hnet30 VSS LPNFET W=0.2U L=0.12U M=1 
X2 net63 net113 VDD VDD LPPFET W=0.62U L=0.12U M=1 
X20 hnet32 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X21 VDD m hnet32 VDD LPPFET W=0.28U L=0.12U M=1 
X22 VDD s net109 VDD LPPFET W=0.62U L=0.12U M=1 
X23 net109 s VSS VSS LPNFET W=0.4U L=0.12U M=1 
X24 VDD s Q VDD LPPFET W=2.4U L=0.12U M=1 
X25 Q s VSS VSS LPNFET W=1.84U L=0.12U M=1 
X26 VDD RN net113 VDD LPPFET W=0.28U L=0.12U M=1 
X27 net113 RN VSS VSS LPNFET W=0.34U L=0.12U M=1 
X28 VDD net100 s VDD LPPFET W=0.66U L=0.12U M=1 
X29 s net100 VSS VSS LPNFET W=0.44U L=0.12U M=1 
X3 net100 SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X30 VDD net109 QN VDD LPPFET W=2.4U L=0.12U M=1 
X31 QN net109 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X32 VDD CKN c VDD LPPFET W=0.44U L=0.12U M=1 
X33 c CKN VSS VSS LPNFET W=0.32U L=0.12U M=1 
X34 VDD c cn VDD LPPFET W=0.28U L=0.12U M=1 
X35 cn c VSS VSS LPNFET W=0.2U L=0.12U M=1 
X4 net73 s net63 VDD LPPFET W=0.28U L=0.12U M=1 
X5 net100 c net73 VDD LPPFET W=0.28U L=0.12U M=1 
X6 net100 cn m VDD LPPFET W=0.3U L=0.12U M=1 
X7 m net113 net94 VSS LPNFET W=0.2U L=0.12U M=1 
X8 m pm net94 VSS LPNFET W=0.34U L=0.12U M=1 
X9 net100 net113 net94 VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS DFFNSRX4TS 

**** 
*.SUBCKT DFFNSRXLTS Q QN CKN D RN SN 
.SUBCKT DFFNSRXLTS Q QN CKN D RN SN VSS VDD
X0 m SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X1 m pm net63 VDD LPPFET W=0.42U L=0.12U M=1 
X10 net91 s net94 VSS LPNFET W=0.2U L=0.12U M=1 
X11 net94 SN VSS VSS LPNFET W=0.4U L=0.12U M=1 
X12 net100 cn net91 VSS LPNFET W=0.2U L=0.12U M=1 
X13 net100 c m VSS LPNFET W=0.2U L=0.12U M=1 
X14 hnet24 D VSS VSS LPNFET W=0.2U L=0.12U M=1 
X15 pm cn hnet24 VSS LPNFET W=0.2U L=0.12U M=1 
X16 hnet26 c pm VDD LPPFET W=0.28U L=0.12U M=1 
X17 VDD D hnet26 VDD LPPFET W=0.28U L=0.12U M=1 
X18 hnet30 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X19 pm c hnet30 VSS LPNFET W=0.2U L=0.12U M=1 
X2 net63 net113 VDD VDD LPPFET W=0.56U L=0.12U M=1 
X20 hnet32 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X21 VDD m hnet32 VDD LPPFET W=0.28U L=0.12U M=1 
X22 VDD s net109 VDD LPPFET W=0.28U L=0.12U M=1 
X23 net109 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X24 VDD s Q VDD LPPFET W=0.34U L=0.12U M=1 
X25 Q s VSS VSS LPNFET W=0.24U L=0.12U M=1 
X26 VDD RN net113 VDD LPPFET W=0.28U L=0.12U M=1 
X27 net113 RN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X28 VDD net100 s VDD LPPFET W=0.28U L=0.12U M=1 
X29 s net100 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 net100 SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X30 VDD net109 QN VDD LPPFET W=0.34U L=0.12U M=1 
X31 QN net109 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X32 VDD CKN c VDD LPPFET W=0.42U L=0.12U M=1 
X33 c CKN VSS VSS LPNFET W=0.3U L=0.12U M=1 
X34 VDD c cn VDD LPPFET W=0.28U L=0.12U M=1 
X35 cn c VSS VSS LPNFET W=0.2U L=0.12U M=1 
X4 net73 s net63 VDD LPPFET W=0.28U L=0.12U M=1 
X5 net100 c net73 VDD LPPFET W=0.28U L=0.12U M=1 
X6 net100 cn m VDD LPPFET W=0.28U L=0.12U M=1 
X7 m net113 net94 VSS LPNFET W=0.2U L=0.12U M=1 
X8 m pm net94 VSS LPNFET W=0.3U L=0.12U M=1 
X9 net100 net113 net94 VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS DFFNSRXLTS 

**** 
*.SUBCKT DFFQX1TS Q CK D 
.SUBCKT DFFQX1TS Q CK D VSS VDD
X0 net37 c m VSS LPNFET W=0.2U L=0.12U M=1 
X1 net37 cn m VDD LPPFET W=0.28U L=0.12U M=1 
X10 hnet29 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X11 pm c hnet29 VSS LPNFET W=0.2U L=0.12U M=1 
X12 hnet31 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X13 VDD m hnet31 VDD LPPFET W=0.28U L=0.12U M=1 
X14 VDD net37 s VDD LPPFET W=0.28U L=0.12U M=1 
X15 s net37 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X16 VDD pm m VDD LPPFET W=0.28U L=0.12U M=1 
X17 m pm VSS VSS LPNFET W=0.2U L=0.12U M=1 
X18 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X19 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 hnet13 D VSS VSS LPNFET W=0.2U L=0.12U M=1 
X20 VDD CK cn VDD LPPFET W=0.38U L=0.12U M=1 
X21 cn CK VSS VSS LPNFET W=0.28U L=0.12U M=1 
X22 VDD s Q VDD LPPFET W=0.64U L=0.12U M=1 
X23 Q s VSS VSS LPNFET W=0.48U L=0.12U M=1 
X3 pm cn hnet13 VSS LPNFET W=0.2U L=0.12U M=1 
X4 hnet15 c pm VDD LPPFET W=0.28U L=0.12U M=1 
X5 VDD D hnet15 VDD LPPFET W=0.28U L=0.12U M=1 
X6 hnet21 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X7 net37 cn hnet21 VSS LPNFET W=0.2U L=0.12U M=1 
X8 hnet23 c net37 VDD LPPFET W=0.28U L=0.12U M=1 
X9 VDD s hnet23 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS DFFQX1TS 

**** 
*.SUBCKT DFFQX2TS Q CK D 
.SUBCKT DFFQX2TS Q CK D VSS VDD
X0 net37 c m VSS LPNFET W=0.2U L=0.12U M=1 
X1 net37 cn m VDD LPPFET W=0.28U L=0.12U M=1 
X10 hnet29 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X11 pm c hnet29 VSS LPNFET W=0.2U L=0.12U M=1 
X12 hnet31 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X13 VDD m hnet31 VDD LPPFET W=0.28U L=0.12U M=1 
X14 VDD net37 s VDD LPPFET W=0.28U L=0.12U M=1 
X15 s net37 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X16 VDD pm m VDD LPPFET W=0.28U L=0.12U M=1 
X17 m pm VSS VSS LPNFET W=0.2U L=0.12U M=1 
X18 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X19 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 hnet13 D VSS VSS LPNFET W=0.2U L=0.12U M=1 
X20 VDD CK cn VDD LPPFET W=0.38U L=0.12U M=1 
X21 cn CK VSS VSS LPNFET W=0.28U L=0.12U M=1 
X22 VDD s Q VDD LPPFET W=1.28U L=0.12U M=1 
X23 Q s VSS VSS LPNFET W=0.92U L=0.12U M=1 
X3 pm cn hnet13 VSS LPNFET W=0.2U L=0.12U M=1 
X4 hnet15 c pm VDD LPPFET W=0.28U L=0.12U M=1 
X5 VDD D hnet15 VDD LPPFET W=0.28U L=0.12U M=1 
X6 hnet21 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X7 net37 cn hnet21 VSS LPNFET W=0.2U L=0.12U M=1 
X8 hnet23 c net37 VDD LPPFET W=0.28U L=0.12U M=1 
X9 VDD s hnet23 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS DFFQX2TS 

**** 
*.SUBCKT DFFQX4TS Q CK D 
.SUBCKT DFFQX4TS Q CK D VSS VDD
X0 net37 c m VSS LPNFET W=0.2U L=0.12U M=1 
X1 net37 cn m VDD LPPFET W=0.28U L=0.12U M=1 
X10 hnet29 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X11 pm c hnet29 VSS LPNFET W=0.2U L=0.12U M=1 
X12 hnet31 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X13 VDD m hnet31 VDD LPPFET W=0.28U L=0.12U M=1 
X14 VDD net37 s VDD LPPFET W=0.5U L=0.12U M=1 
X15 s net37 VSS VSS LPNFET W=0.36U L=0.12U M=1 
X16 VDD pm m VDD LPPFET W=0.28U L=0.12U M=1 
X17 m pm VSS VSS LPNFET W=0.2U L=0.12U M=1 
X18 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X19 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 hnet13 D VSS VSS LPNFET W=0.2U L=0.12U M=1 
X20 VDD CK cn VDD LPPFET W=0.38U L=0.12U M=1 
X21 cn CK VSS VSS LPNFET W=0.28U L=0.12U M=1 
X22 VDD s Q VDD LPPFET W=2.56U L=0.12U M=1 
X23 Q s VSS VSS LPNFET W=1.74U L=0.12U M=1 
X3 pm cn hnet13 VSS LPNFET W=0.2U L=0.12U M=1 
X4 hnet15 c pm VDD LPPFET W=0.28U L=0.12U M=1 
X5 VDD D hnet15 VDD LPPFET W=0.28U L=0.12U M=1 
X6 hnet21 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X7 net37 cn hnet21 VSS LPNFET W=0.2U L=0.12U M=1 
X8 hnet23 c net37 VDD LPPFET W=0.28U L=0.12U M=1 
X9 VDD s hnet23 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS DFFQX4TS 

**** 
*.SUBCKT DFFQXLTS Q CK D 
.SUBCKT DFFQXLTS Q CK D VSS VDD
X0 net37 c m VSS LPNFET W=0.2U L=0.12U M=1 
X1 net37 cn m VDD LPPFET W=0.28U L=0.12U M=1 
X10 hnet29 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X11 pm c hnet29 VSS LPNFET W=0.2U L=0.12U M=1 
X12 hnet31 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X13 VDD m hnet31 VDD LPPFET W=0.28U L=0.12U M=1 
X14 VDD net37 s VDD LPPFET W=0.28U L=0.12U M=1 
X15 s net37 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X16 VDD pm m VDD LPPFET W=0.28U L=0.12U M=1 
X17 m pm VSS VSS LPNFET W=0.2U L=0.12U M=1 
X18 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X19 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 hnet13 D VSS VSS LPNFET W=0.2U L=0.12U M=1 
X20 VDD CK cn VDD LPPFET W=0.38U L=0.12U M=1 
X21 cn CK VSS VSS LPNFET W=0.28U L=0.12U M=1 
X22 VDD s Q VDD LPPFET W=0.34U L=0.12U M=1 
X23 Q s VSS VSS LPNFET W=0.24U L=0.12U M=1 
X3 pm cn hnet13 VSS LPNFET W=0.2U L=0.12U M=1 
X4 hnet15 c pm VDD LPPFET W=0.28U L=0.12U M=1 
X5 VDD D hnet15 VDD LPPFET W=0.28U L=0.12U M=1 
X6 hnet21 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X7 net37 cn hnet21 VSS LPNFET W=0.2U L=0.12U M=1 
X8 hnet23 c net37 VDD LPPFET W=0.28U L=0.12U M=1 
X9 VDD s hnet23 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS DFFQXLTS 

**** 
*.SUBCKT DFFRHQX1TS Q CK D RN 
.SUBCKT DFFRHQX1TS Q CK D RN VSS VDD
X0 VDD c hnet24 VDD LPPFET W=0.6U L=0.12U M=1 
X1 hnet24 nmin pm VDD LPPFET W=0.6U L=0.12U M=1 
X10 net81 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X11 m RN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X12 m pm VDD VDD LPPFET W=0.96U L=0.12U M=1 
X13 net105 cn m VDD LPPFET W=0.92U L=0.12U M=1 
X14 cn CK VSS VSS LPNFET W=0.2U L=0.12U M=1 
X15 net98 RN net102 VSS LPNFET W=0.2U L=0.12U M=1 
X16 net105 cn net98 VSS LPNFET W=0.2U L=0.12U M=1 
X17 net102 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X18 net105 c m VSS LPNFET W=0.48U L=0.12U M=1 
X19 hnet34 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 hnet28 cn VSS VSS LPNFET W=0.44U L=0.12U M=1 
X20 pm c hnet34 VSS LPNFET W=0.2U L=0.12U M=1 
X21 hnet36 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X22 VDD m hnet36 VDD LPPFET W=0.28U L=0.12U M=1 
X23 VDD D nmin VDD LPPFET W=0.28U L=0.12U M=1 
X24 nmin D VSS VSS LPNFET W=0.2U L=0.12U M=1 
X25 VDD net105 s VDD LPPFET W=0.28U L=0.12U M=1 
X26 s net105 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X27 VDD net105 Q VDD LPPFET W=0.74U L=0.12U M=1 
X28 Q net105 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X29 VDD net118 c VDD LPPFET W=0.84U L=0.12U M=1 
X3 pm nmin hnet28 VSS LPNFET W=0.44U L=0.12U M=1 
X30 c net118 VSS VSS LPNFET W=0.3U L=0.12U M=1 
X31 VDD CK net118 VDD LPPFET W=0.28U L=0.12U M=1 
X32 net118 CK VSS VSS LPNFET W=0.28U L=0.12U M=1 
X4 hnet32 RN VSS VSS LPNFET W=0.58U L=0.12U M=1 
X5 m pm hnet32 VSS LPNFET W=0.58U L=0.12U M=1 
X6 net71 CK VDD VDD LPPFET W=0.7U L=0.12U M=1 
X7 cn c net71 VDD LPPFET W=0.52U L=0.12U M=1 
X8 net105 RN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X9 net105 c net81 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS DFFRHQX1TS 

**** 
*.SUBCKT DFFRHQX2TS Q CK D RN 
.SUBCKT DFFRHQX2TS Q CK D RN VSS VDD
X0 VDD c hnet24 VDD LPPFET W=1.02U L=0.12U M=1 
X1 hnet24 nmin pm VDD LPPFET W=1.02U L=0.12U M=1 
X10 net77 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X11 m RN VDD VDD LPPFET W=0.4U L=0.12U M=1 
X12 m pm VDD VDD LPPFET W=1.6U L=0.12U M=1 
X13 net105 cn m VDD LPPFET W=1.54U L=0.12U M=1 
X14 cn CK VSS VSS LPNFET W=0.28U L=0.12U M=1 
X15 net98 RN net95 VSS LPNFET W=0.2U L=0.12U M=1 
X16 net105 cn net98 VSS LPNFET W=0.2U L=0.12U M=1 
X17 net95 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X18 net105 c m VSS LPNFET W=0.66U L=0.12U M=1 
X19 hnet34 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 hnet28 cn VSS VSS LPNFET W=0.74U L=0.12U M=1 
X20 pm c hnet34 VSS LPNFET W=0.2U L=0.12U M=1 
X21 hnet36 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X22 VDD m hnet36 VDD LPPFET W=0.28U L=0.12U M=1 
X23 VDD D nmin VDD LPPFET W=0.36U L=0.12U M=1 
X24 nmin D VSS VSS LPNFET W=0.28U L=0.12U M=1 
X25 VDD net105 s VDD LPPFET W=0.28U L=0.12U M=1 
X26 s net105 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X27 VDD net105 Q VDD LPPFET W=1.3U L=0.12U M=1 
X28 Q net105 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X29 VDD net118 c VDD LPPFET W=1.16U L=0.12U M=1 
X3 pm nmin hnet28 VSS LPNFET W=0.74U L=0.12U M=1 
X30 c net118 VSS VSS LPNFET W=0.44U L=0.12U M=1 
X31 VDD CK net118 VDD LPPFET W=0.34U L=0.12U M=1 
X32 net118 CK VSS VSS LPNFET W=0.34U L=0.12U M=1 
X4 hnet32 RN VSS VSS LPNFET W=0.98U L=0.12U M=1 
X5 m pm hnet32 VSS LPNFET W=0.98U L=0.12U M=1 
X6 net71 CK VDD VDD LPPFET W=0.98U L=0.12U M=1 
X7 cn c net71 VDD LPPFET W=0.74U L=0.12U M=1 
X8 net105 RN VDD VDD LPPFET W=0.4U L=0.12U M=1 
X9 net105 c net77 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS DFFRHQX2TS 

**** 
*.SUBCKT DFFRHQX4TS Q CK D RN 
.SUBCKT DFFRHQX4TS Q CK D RN VSS VDD
X0 VDD c hnet25 VDD LPPFET W=0.96U L=0.12U M=1 
X1 hnet25 nmin pm VDD LPPFET W=0.96U L=0.12U M=1 
X10 hnet31 RN VSS VSS LPNFET W=0.82U L=0.12U M=1 
X11 m pm hnet31 VSS LPNFET W=0.82U L=0.12U M=1 
X12 net71 CK VDD VDD LPPFET W=1.3U L=0.12U M=1 
X13 cn c net71 VDD LPPFET W=1.26U L=0.12U M=1 
X14 net105 RN VDD VDD LPPFET W=0.7U L=0.12U M=1 
X15 net105 c net77 VDD LPPFET W=0.28U L=0.12U M=1 
X16 net77 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X17 m RN VDD VDD LPPFET W=0.7U L=0.12U M=1 
X18 m pm VDD VDD LPPFET W=2.56U L=0.12U M=1 
X19 net105 cn m VDD LPPFET W=2.8U L=0.12U M=1 
X2 VDD c hnet22 VDD LPPFET W=0.96U L=0.12U M=1 
X20 cn CK VSS VSS LPNFET W=0.48U L=0.12U M=1 
X21 net98 RN net95 VSS LPNFET W=0.2U L=0.12U M=1 
X22 net105 cn net98 VSS LPNFET W=0.2U L=0.12U M=1 
X23 net95 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X24 net105 c m VSS LPNFET W=1.48U L=0.12U M=1 
X25 hnet37 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X26 pm c hnet37 VSS LPNFET W=0.2U L=0.12U M=1 
X27 hnet39 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X28 VDD m hnet39 VDD LPPFET W=0.28U L=0.12U M=1 
X29 VDD D nmin VDD LPPFET W=0.66U L=0.12U M=1 
X3 hnet22 nmin pm VDD LPPFET W=0.96U L=0.12U M=1 
X30 nmin D VSS VSS LPNFET W=0.48U L=0.12U M=1 
X31 VDD net105 s VDD LPPFET W=0.28U L=0.12U M=1 
X32 s net105 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X33 VDD net105 Q VDD LPPFET W=2.6U L=0.12U M=1 
X34 Q net105 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X35 VDD net118 c VDD LPPFET W=2.06U L=0.12U M=1 
X36 c net118 VSS VSS LPNFET W=0.74U L=0.12U M=1 
X37 VDD CK net118 VDD LPPFET W=0.56U L=0.12U M=1 
X38 net118 CK VSS VSS LPNFET W=0.56U L=0.12U M=1 
X4 hnet30 cn VSS VSS LPNFET W=0.7U L=0.12U M=1 
X5 pm nmin hnet30 VSS LPNFET W=0.7U L=0.12U M=1 
X6 hnet26 cn VSS VSS LPNFET W=0.7U L=0.12U M=1 
X7 pm nmin hnet26 VSS LPNFET W=0.7U L=0.12U M=1 
X8 hnet35 RN VSS VSS LPNFET W=0.82U L=0.12U M=1 
X9 m pm hnet35 VSS LPNFET W=0.82U L=0.12U M=1 
.ENDS DFFRHQX4TS 

**** 
*.SUBCKT DFFRHQX8TS Q CK D RN 
.SUBCKT DFFRHQX8TS Q CK D RN VSS VDD
X0 VDD c hnet25 VDD LPPFET W=0.96U L=0.12U M=1 
X1 hnet25 nmin pm VDD LPPFET W=0.96U L=0.12U M=1 
X10 hnet31 RN VSS VSS LPNFET W=0.82U L=0.12U M=1 
X11 m pm hnet31 VSS LPNFET W=0.82U L=0.12U M=1 
X12 net71 CK VDD VDD LPPFET W=1.3U L=0.12U M=1 
X13 cn c net71 VDD LPPFET W=1.26U L=0.12U M=1 
X14 net105 RN VDD VDD LPPFET W=0.7U L=0.12U M=1 
X15 net105 c net81 VDD LPPFET W=0.28U L=0.12U M=1 
X16 net81 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X17 m RN VDD VDD LPPFET W=0.7U L=0.12U M=1 
X18 m pm VDD VDD LPPFET W=2.56U L=0.12U M=1 
X19 net105 cn m VDD LPPFET W=2.8U L=0.12U M=1 
X2 VDD c hnet22 VDD LPPFET W=0.96U L=0.12U M=1 
X20 cn CK VSS VSS LPNFET W=0.48U L=0.12U M=1 
X21 net98 RN net102 VSS LPNFET W=0.2U L=0.12U M=1 
X22 net105 cn net98 VSS LPNFET W=0.2U L=0.12U M=1 
X23 net102 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X24 net105 c m VSS LPNFET W=1.48U L=0.12U M=1 
X25 hnet37 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X26 pm c hnet37 VSS LPNFET W=0.2U L=0.12U M=1 
X27 hnet39 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X28 VDD m hnet39 VDD LPPFET W=0.28U L=0.12U M=1 
X29 VDD D nmin VDD LPPFET W=0.66U L=0.12U M=1 
X3 hnet22 nmin pm VDD LPPFET W=0.96U L=0.12U M=1 
X30 nmin D VSS VSS LPNFET W=0.48U L=0.12U M=1 
X31 VDD net105 s VDD LPPFET W=0.28U L=0.12U M=1 
X32 s net105 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X33 VDD net105 Q VDD LPPFET W=5.2U L=0.12U M=1 
X34 Q net105 VSS VSS LPNFET W=3.68U L=0.12U M=1 
X35 VDD net118 c VDD LPPFET W=2.06U L=0.12U M=1 
X36 c net118 VSS VSS LPNFET W=0.74U L=0.12U M=1 
X37 VDD CK net118 VDD LPPFET W=0.56U L=0.12U M=1 
X38 net118 CK VSS VSS LPNFET W=0.56U L=0.12U M=1 
X4 hnet30 cn VSS VSS LPNFET W=0.7U L=0.12U M=1 
X5 pm nmin hnet30 VSS LPNFET W=0.7U L=0.12U M=1 
X6 hnet26 cn VSS VSS LPNFET W=0.7U L=0.12U M=1 
X7 pm nmin hnet26 VSS LPNFET W=0.7U L=0.12U M=1 
X8 hnet35 RN VSS VSS LPNFET W=0.82U L=0.12U M=1 
X9 m pm hnet35 VSS LPNFET W=0.82U L=0.12U M=1 
.ENDS DFFRHQX8TS 

**** 
*.SUBCKT DFFRX1TS Q QN CK D RN 
.SUBCKT DFFRX1TS Q QN CK D RN VSS VDD
X0 hnet22 RN VSS VSS LPNFET W=0.32U L=0.12U M=1 
X1 s net88 hnet22 VSS LPNFET W=0.32U L=0.12U M=1 
X10 pm c hnet31 VSS LPNFET W=0.2U L=0.12U M=1 
X11 hnet42 RN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X12 hnet37 D hnet42 VSS LPNFET W=0.2U L=0.12U M=1 
X13 pm cn hnet37 VSS LPNFET W=0.2U L=0.12U M=1 
X14 pm RN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X15 net88 c net72 VDD LPPFET W=0.28U L=0.12U M=1 
X16 net72 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X17 net88 cn m VDD LPPFET W=0.28U L=0.12U M=1 
X18 net88 cn net85 VSS LPNFET W=0.2U L=0.12U M=1 
X19 net85 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 VDD RN s VDD LPPFET W=0.28U L=0.12U M=1 
X20 net88 c m VSS LPNFET W=0.2U L=0.12U M=1 
X21 VDD s net89 VDD LPPFET W=0.28U L=0.12U M=1 
X22 net89 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X23 VDD pm m VDD LPPFET W=0.28U L=0.12U M=1 
X24 m pm VSS VSS LPNFET W=0.2U L=0.12U M=1 
X25 VDD s Q VDD LPPFET W=0.64U L=0.12U M=1 
X26 Q s VSS VSS LPNFET W=0.46U L=0.12U M=1 
X27 VDD net89 QN VDD LPPFET W=0.64U L=0.12U M=1 
X28 QN net89 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X29 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X3 VDD net88 s VDD LPPFET W=0.28U L=0.12U M=1 
X30 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X31 VDD CK cn VDD LPPFET W=0.42U L=0.12U M=1 
X32 cn CK VSS VSS LPNFET W=0.3U L=0.12U M=1 
X4 VDD m hnet26 VDD LPPFET W=0.28U L=0.12U M=1 
X5 hnet26 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X6 VDD D hnet30 VDD LPPFET W=0.28U L=0.12U M=1 
X7 hnet30 c pm VDD LPPFET W=0.28U L=0.12U M=1 
X8 hnet36 RN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X9 hnet31 m hnet36 VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS DFFRX1TS 

**** 
*.SUBCKT DFFRX2TS Q QN CK D RN 
.SUBCKT DFFRX2TS Q QN CK D RN VSS VDD
X0 hnet22 RN VSS VSS LPNFET W=0.52U L=0.12U M=1 
X1 s net88 hnet22 VSS LPNFET W=0.52U L=0.12U M=1 
X10 pm c hnet31 VSS LPNFET W=0.2U L=0.12U M=1 
X11 hnet42 RN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X12 hnet37 D hnet42 VSS LPNFET W=0.2U L=0.12U M=1 
X13 pm cn hnet37 VSS LPNFET W=0.2U L=0.12U M=1 
X14 pm RN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X15 net88 c net72 VDD LPPFET W=0.28U L=0.12U M=1 
X16 net72 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X17 net88 cn m VDD LPPFET W=0.28U L=0.12U M=1 
X18 net88 cn net85 VSS LPNFET W=0.2U L=0.12U M=1 
X19 net85 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 VDD RN s VDD LPPFET W=0.38U L=0.12U M=1 
X20 net88 c m VSS LPNFET W=0.2U L=0.12U M=1 
X21 VDD s net89 VDD LPPFET W=0.3U L=0.12U M=1 
X22 net89 s VSS VSS LPNFET W=0.22U L=0.12U M=1 
X23 VDD pm m VDD LPPFET W=0.28U L=0.12U M=1 
X24 m pm VSS VSS LPNFET W=0.2U L=0.12U M=1 
X25 VDD s Q VDD LPPFET W=1.28U L=0.12U M=1 
X26 Q s VSS VSS LPNFET W=0.92U L=0.12U M=1 
X27 VDD net89 QN VDD LPPFET W=1.28U L=0.12U M=1 
X28 QN net89 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X29 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X3 VDD net88 s VDD LPPFET W=0.38U L=0.12U M=1 
X30 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X31 VDD CK cn VDD LPPFET W=0.42U L=0.12U M=1 
X32 cn CK VSS VSS LPNFET W=0.3U L=0.12U M=1 
X4 VDD m hnet26 VDD LPPFET W=0.28U L=0.12U M=1 
X5 hnet26 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X6 VDD D hnet30 VDD LPPFET W=0.28U L=0.12U M=1 
X7 hnet30 c pm VDD LPPFET W=0.28U L=0.12U M=1 
X8 hnet36 RN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X9 hnet31 m hnet36 VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS DFFRX2TS 

**** 
*.SUBCKT DFFRX4TS Q QN CK D RN 
.SUBCKT DFFRX4TS Q QN CK D RN VSS VDD
X0 hnet22 RN VSS VSS LPNFET W=0.92U L=0.12U M=1 
X1 s net88 hnet22 VSS LPNFET W=0.92U L=0.12U M=1 
X10 pm c hnet31 VSS LPNFET W=0.2U L=0.12U M=1 
X11 hnet42 RN VSS VSS LPNFET W=0.24U L=0.12U M=1 
X12 hnet37 D hnet42 VSS LPNFET W=0.24U L=0.12U M=1 
X13 pm cn hnet37 VSS LPNFET W=0.24U L=0.12U M=1 
X14 pm RN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X15 net88 c net72 VDD LPPFET W=0.28U L=0.12U M=1 
X16 net72 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X17 net88 cn m VDD LPPFET W=0.48U L=0.12U M=1 
X18 net88 cn net85 VSS LPNFET W=0.2U L=0.12U M=1 
X19 net85 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 VDD RN s VDD LPPFET W=0.62U L=0.12U M=1 
X20 net88 c m VSS LPNFET W=0.34U L=0.12U M=1 
X21 VDD s net89 VDD LPPFET W=0.62U L=0.12U M=1 
X22 net89 s VSS VSS LPNFET W=0.44U L=0.12U M=1 
X23 VDD pm m VDD LPPFET W=0.48U L=0.12U M=1 
X24 m pm VSS VSS LPNFET W=0.34U L=0.12U M=1 
X25 VDD s Q VDD LPPFET W=2.56U L=0.12U M=1 
X26 Q s VSS VSS LPNFET W=1.84U L=0.12U M=1 
X27 VDD net89 QN VDD LPPFET W=2.56U L=0.12U M=1 
X28 QN net89 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X29 VDD cn c VDD LPPFET W=0.34U L=0.12U M=1 
X3 VDD net88 s VDD LPPFET W=0.62U L=0.12U M=1 
X30 c cn VSS VSS LPNFET W=0.24U L=0.12U M=1 
X31 VDD CK cn VDD LPPFET W=0.52U L=0.12U M=1 
X32 cn CK VSS VSS LPNFET W=0.38U L=0.12U M=1 
X4 VDD m hnet26 VDD LPPFET W=0.28U L=0.12U M=1 
X5 hnet26 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X6 VDD D hnet30 VDD LPPFET W=0.28U L=0.12U M=1 
X7 hnet30 c pm VDD LPPFET W=0.28U L=0.12U M=1 
X8 hnet36 RN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X9 hnet31 m hnet36 VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS DFFRX4TS 

**** 
*.SUBCKT DFFRXLTS Q QN CK D RN 
.SUBCKT DFFRXLTS Q QN CK D RN VSS VDD
X0 hnet22 RN VSS VSS LPNFET W=0.22U L=0.12U M=1 
X1 s net88 hnet22 VSS LPNFET W=0.22U L=0.12U M=1 
X10 pm c hnet31 VSS LPNFET W=0.2U L=0.12U M=1 
X11 hnet42 RN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X12 hnet37 D hnet42 VSS LPNFET W=0.2U L=0.12U M=1 
X13 pm cn hnet37 VSS LPNFET W=0.2U L=0.12U M=1 
X14 pm RN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X15 net88 c net72 VDD LPPFET W=0.28U L=0.12U M=1 
X16 net72 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X17 net88 cn m VDD LPPFET W=0.28U L=0.12U M=1 
X18 net88 cn net85 VSS LPNFET W=0.2U L=0.12U M=1 
X19 net85 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 VDD RN s VDD LPPFET W=0.28U L=0.12U M=1 
X20 net88 c m VSS LPNFET W=0.2U L=0.12U M=1 
X21 VDD s net89 VDD LPPFET W=0.28U L=0.12U M=1 
X22 net89 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X23 VDD pm m VDD LPPFET W=0.28U L=0.12U M=1 
X24 m pm VSS VSS LPNFET W=0.2U L=0.12U M=1 
X25 VDD s Q VDD LPPFET W=0.34U L=0.12U M=1 
X26 Q s VSS VSS LPNFET W=0.24U L=0.12U M=1 
X27 VDD net89 QN VDD LPPFET W=0.34U L=0.12U M=1 
X28 QN net89 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X29 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X3 VDD net88 s VDD LPPFET W=0.28U L=0.12U M=1 
X30 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X31 VDD CK cn VDD LPPFET W=0.42U L=0.12U M=1 
X32 cn CK VSS VSS LPNFET W=0.3U L=0.12U M=1 
X4 VDD m hnet26 VDD LPPFET W=0.28U L=0.12U M=1 
X5 hnet26 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X6 VDD D hnet30 VDD LPPFET W=0.28U L=0.12U M=1 
X7 hnet30 c pm VDD LPPFET W=0.28U L=0.12U M=1 
X8 hnet36 RN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X9 hnet31 m hnet36 VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS DFFRXLTS 

**** 
*.SUBCKT DFFSHQX1TS Q CK D SN 
.SUBCKT DFFSHQX1TS Q CK D SN VSS VDD
X0 VDD c hnet25 VDD LPPFET W=0.52U L=0.12U M=1 
X1 hnet25 nmin pm VDD LPPFET W=0.52U L=0.12U M=1 
X10 net76 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X11 net94 cn m VDD LPPFET W=0.96U L=0.12U M=1 
X12 cn CK VSS VSS LPNFET W=0.2U L=0.12U M=1 
X13 net94 cn net88 VSS LPNFET W=0.2U L=0.12U M=1 
X14 net88 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X15 net94 nmset VSS VSS LPNFET W=0.2U L=0.12U M=1 
X16 net94 c m VSS LPNFET W=0.48U L=0.12U M=1 
X17 hnet33 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X18 pm c hnet33 VSS LPNFET W=0.2U L=0.12U M=1 
X19 hnet35 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X2 hnet31 SN VSS VSS LPNFET W=0.56U L=0.12U M=1 
X20 VDD m hnet35 VDD LPPFET W=0.28U L=0.12U M=1 
X21 VDD pm m VDD LPPFET W=0.96U L=0.12U M=1 
X22 m pm VSS VSS LPNFET W=0.5U L=0.12U M=1 
X23 VDD SN nmset VDD LPPFET W=0.28U L=0.12U M=1 
X24 nmset SN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X25 VDD D nmin VDD LPPFET W=0.28U L=0.12U M=1 
X26 nmin D VSS VSS LPNFET W=0.2U L=0.12U M=1 
X27 VDD net94 s VDD LPPFET W=0.28U L=0.12U M=1 
X28 s net94 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X29 VDD net94 Q VDD LPPFET W=0.74U L=0.12U M=1 
X3 hnet26 cn hnet31 VSS LPNFET W=0.56U L=0.12U M=1 
X30 Q net94 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X31 VDD net111 c VDD LPPFET W=0.72U L=0.12U M=1 
X32 c net111 VSS VSS LPNFET W=0.26U L=0.12U M=1 
X33 VDD CK net111 VDD LPPFET W=0.28U L=0.12U M=1 
X34 net111 CK VSS VSS LPNFET W=0.28U L=0.12U M=1 
X4 pm nmin hnet26 VSS LPNFET W=0.56U L=0.12U M=1 
X5 net61 CK VDD VDD LPPFET W=0.62U L=0.12U M=1 
X6 cn c net61 VDD LPPFET W=0.52U L=0.12U M=1 
X7 pm SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X8 net70 nmset net76 VDD LPPFET W=0.28U L=0.12U M=1 
X9 net94 c net70 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS DFFSHQX1TS 

**** 
*.SUBCKT DFFSHQX2TS Q CK D SN 
.SUBCKT DFFSHQX2TS Q CK D SN VSS VDD
X0 VDD c hnet25 VDD LPPFET W=0.9U L=0.12U M=1 
X1 hnet25 nmin pm VDD LPPFET W=0.9U L=0.12U M=1 
X10 net76 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X11 net94 cn m VDD LPPFET W=1.64U L=0.12U M=1 
X12 cn CK VSS VSS LPNFET W=0.3U L=0.12U M=1 
X13 net94 cn net88 VSS LPNFET W=0.2U L=0.12U M=1 
X14 net88 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X15 net94 nmset VSS VSS LPNFET W=0.28U L=0.12U M=1 
X16 net94 c m VSS LPNFET W=0.82U L=0.12U M=1 
X17 hnet33 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X18 pm c hnet33 VSS LPNFET W=0.2U L=0.12U M=1 
X19 hnet35 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X2 hnet31 SN VSS VSS LPNFET W=0.9U L=0.12U M=1 
X20 VDD m hnet35 VDD LPPFET W=0.28U L=0.12U M=1 
X21 VDD pm m VDD LPPFET W=1.64U L=0.12U M=1 
X22 m pm VSS VSS LPNFET W=0.86U L=0.12U M=1 
X23 VDD SN nmset VDD LPPFET W=0.28U L=0.12U M=1 
X24 nmset SN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X25 VDD D nmin VDD LPPFET W=0.36U L=0.12U M=1 
X26 nmin D VSS VSS LPNFET W=0.28U L=0.12U M=1 
X27 VDD net94 s VDD LPPFET W=0.28U L=0.12U M=1 
X28 s net94 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X29 VDD net94 Q VDD LPPFET W=1.48U L=0.12U M=1 
X3 hnet26 cn hnet31 VSS LPNFET W=0.9U L=0.12U M=1 
X30 Q net94 VSS VSS LPNFET W=0.84U L=0.12U M=1 
X31 VDD net111 c VDD LPPFET W=1.16U L=0.12U M=1 
X32 c net111 VSS VSS LPNFET W=0.42U L=0.12U M=1 
X33 VDD CK net111 VDD LPPFET W=0.32U L=0.12U M=1 
X34 net111 CK VSS VSS LPNFET W=0.32U L=0.12U M=1 
X4 pm nmin hnet26 VSS LPNFET W=0.9U L=0.12U M=1 
X5 net63 CK VDD VDD LPPFET W=1.06U L=0.12U M=1 
X6 cn c net63 VDD LPPFET W=0.8U L=0.12U M=1 
X7 pm SN VDD VDD LPPFET W=0.34U L=0.12U M=1 
X8 net72 nmset net76 VDD LPPFET W=0.28U L=0.12U M=1 
X9 net94 c net72 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS DFFSHQX2TS 

**** 
*.SUBCKT DFFSHQX4TS Q CK D SN 
.SUBCKT DFFSHQX4TS Q CK D SN VSS VDD
X0 hnet28 SN VSS VSS LPNFET W=0.76U L=0.12U M=1 
X1 hnet22 cn hnet28 VSS LPNFET W=0.76U L=0.12U M=1 
X10 net63 CK VDD VDD LPPFET W=1.84U L=0.12U M=1 
X11 cn c net63 VDD LPPFET W=1.3U L=0.12U M=1 
X12 pm SN VDD VDD LPPFET W=0.64U L=0.12U M=1 
X13 net72 nmset net76 VDD LPPFET W=0.28U L=0.12U M=1 
X14 net94 c net72 VDD LPPFET W=0.28U L=0.12U M=1 
X15 net76 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X16 net94 cn m VDD LPPFET W=2.38U L=0.12U M=1 
X17 cn CK VSS VSS LPNFET W=0.52U L=0.12U M=1 
X18 net94 cn net88 VSS LPNFET W=0.2U L=0.12U M=1 
X19 net88 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 pm nmin hnet22 VSS LPNFET W=0.76U L=0.12U M=1 
X20 net94 nmset VSS VSS LPNFET W=0.52U L=0.12U M=1 
X21 net94 c m VSS LPNFET W=1.3U L=0.12U M=1 
X22 hnet36 m VSS VSS LPNFET W=0.22U L=0.12U M=1 
X23 pm c hnet36 VSS LPNFET W=0.22U L=0.12U M=1 
X24 hnet38 cn pm VDD LPPFET W=0.3U L=0.12U M=1 
X25 VDD m hnet38 VDD LPPFET W=0.3U L=0.12U M=1 
X26 VDD pm m VDD LPPFET W=2.5U L=0.12U M=1 
X27 m pm VSS VSS LPNFET W=1.3U L=0.12U M=1 
X28 VDD SN nmset VDD LPPFET W=0.28U L=0.12U M=1 
X29 nmset SN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 hnet29 SN VSS VSS LPNFET W=0.76U L=0.12U M=1 
X30 VDD D nmin VDD LPPFET W=0.66U L=0.12U M=1 
X31 nmin D VSS VSS LPNFET W=0.48U L=0.12U M=1 
X32 VDD net94 s VDD LPPFET W=0.28U L=0.12U M=1 
X33 s net94 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X34 VDD net94 Q VDD LPPFET W=2.6U L=0.12U M=1 
X35 Q net94 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X36 VDD net111 c VDD LPPFET W=2.02U L=0.12U M=1 
X37 c net111 VSS VSS LPNFET W=0.72U L=0.12U M=1 
X38 VDD CK net111 VDD LPPFET W=0.54U L=0.12U M=1 
X39 net111 CK VSS VSS LPNFET W=0.54U L=0.12U M=1 
X4 hnet24 cn hnet29 VSS LPNFET W=0.76U L=0.12U M=1 
X5 pm nmin hnet24 VSS LPNFET W=0.76U L=0.12U M=1 
X6 VDD c hnet34 VDD LPPFET W=0.76U L=0.12U M=1 
X7 hnet34 nmin pm VDD LPPFET W=0.76U L=0.12U M=1 
X8 VDD c hnet31 VDD LPPFET W=0.76U L=0.12U M=1 
X9 hnet31 nmin pm VDD LPPFET W=0.76U L=0.12U M=1 
.ENDS DFFSHQX4TS 

**** 
*.SUBCKT DFFSHQX8TS Q CK D SN 
.SUBCKT DFFSHQX8TS Q CK D SN VSS VDD
X0 hnet28 SN VSS VSS LPNFET W=0.8U L=0.12U M=1 
X1 hnet22 cn hnet28 VSS LPNFET W=0.8U L=0.12U M=1 
X10 net61 CK VDD VDD LPPFET W=1.84U L=0.12U M=1 
X11 cn c net61 VDD LPPFET W=1.32U L=0.12U M=1 
X12 pm SN VDD VDD LPPFET W=0.64U L=0.12U M=1 
X13 net70 nmset net76 VDD LPPFET W=0.28U L=0.12U M=1 
X14 net94 c net70 VDD LPPFET W=0.28U L=0.12U M=1 
X15 net76 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X16 net94 cn m VDD LPPFET W=2.66U L=0.12U M=1 
X17 cn CK VSS VSS LPNFET W=0.52U L=0.12U M=1 
X18 net94 cn net88 VSS LPNFET W=0.2U L=0.12U M=1 
X19 net88 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 pm nmin hnet22 VSS LPNFET W=0.8U L=0.12U M=1 
X20 net94 nmset VSS VSS LPNFET W=0.52U L=0.12U M=1 
X21 net94 c m VSS LPNFET W=1.5U L=0.12U M=1 
X22 hnet36 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X23 pm c hnet36 VSS LPNFET W=0.2U L=0.12U M=1 
X24 hnet38 cn pm VDD LPPFET W=0.3U L=0.12U M=1 
X25 VDD m hnet38 VDD LPPFET W=0.3U L=0.12U M=1 
X26 VDD pm m VDD LPPFET W=2.66U L=0.12U M=1 
X27 m pm VSS VSS LPNFET W=1.5U L=0.12U M=1 
X28 VDD SN nmset VDD LPPFET W=0.28U L=0.12U M=1 
X29 nmset SN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 hnet29 SN VSS VSS LPNFET W=0.8U L=0.12U M=1 
X30 VDD D nmin VDD LPPFET W=0.66U L=0.12U M=1 
X31 nmin D VSS VSS LPNFET W=0.48U L=0.12U M=1 
X32 VDD net94 s VDD LPPFET W=0.28U L=0.12U M=1 
X33 s net94 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X34 VDD net94 Q VDD LPPFET W=5.34U L=0.12U M=1 
X35 Q net94 VSS VSS LPNFET W=3.48U L=0.12U M=1 
X36 VDD net111 c VDD LPPFET W=1.98U L=0.12U M=1 
X37 c net111 VSS VSS LPNFET W=0.72U L=0.12U M=1 
X38 VDD CK net111 VDD LPPFET W=0.54U L=0.12U M=1 
X39 net111 CK VSS VSS LPNFET W=0.54U L=0.12U M=1 
X4 hnet24 cn hnet29 VSS LPNFET W=0.8U L=0.12U M=1 
X5 pm nmin hnet24 VSS LPNFET W=0.8U L=0.12U M=1 
X6 VDD c hnet34 VDD LPPFET W=0.82U L=0.12U M=1 
X7 hnet34 nmin pm VDD LPPFET W=0.82U L=0.12U M=1 
X8 VDD c hnet31 VDD LPPFET W=0.82U L=0.12U M=1 
X9 hnet31 nmin pm VDD LPPFET W=0.82U L=0.12U M=1 
.ENDS DFFSHQX8TS 

**** 
*.SUBCKT DFFSRHQX1TS Q CK D RN SN 
.SUBCKT DFFSRHQX1TS Q CK D RN SN VSS VDD
X0 hnet29 SN VSS VSS LPNFET W=0.54U L=0.12U M=1 
X1 hnet24 cn hnet29 VSS LPNFET W=0.54U L=0.12U M=1 
X10 hnet45 nmset net130 VDD LPPFET W=0.26U L=0.12U M=1 
X11 net88 CK VDD VDD LPPFET W=0.7U L=0.12U M=1 
X12 cn c net88 VDD LPPFET W=0.52U L=0.12U M=1 
X13 pm SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X14 m pm VDD VDD LPPFET W=0.66U L=0.12U M=1 
X15 net102 nmset net106 VDD LPPFET W=0.28U L=0.12U M=1 
X16 net130 c net102 VDD LPPFET W=0.28U L=0.12U M=1 
X17 net106 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X18 net130 cn m VDD LPPFET W=0.66U L=0.12U M=1 
X19 cn CK VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 pm nmin hnet24 VSS LPNFET W=0.54U L=0.12U M=1 
X20 net115 RN net114 VSS LPNFET W=0.2U L=0.12U M=1 
X21 net130 cn net115 VSS LPNFET W=0.2U L=0.12U M=1 
X22 net114 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X23 net130 nmset VSS VSS LPNFET W=0.2U L=0.12U M=1 
X24 m nmset VSS VSS LPNFET W=0.2U L=0.12U M=1 
X25 net130 c m VSS LPNFET W=0.48U L=0.12U M=1 
X26 hnet47 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X27 pm c hnet47 VSS LPNFET W=0.2U L=0.12U M=1 
X28 hnet49 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X29 VDD m hnet49 VDD LPPFET W=0.28U L=0.12U M=1 
X3 hnet33 RN VSS VSS LPNFET W=0.5U L=0.12U M=1 
X30 VDD SN nmset VDD LPPFET W=0.28U L=0.12U M=1 
X31 nmset SN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X32 VDD D nmin VDD LPPFET W=0.28U L=0.12U M=1 
X33 nmin D VSS VSS LPNFET W=0.2U L=0.12U M=1 
X34 VDD net130 s VDD LPPFET W=0.28U L=0.12U M=1 
X35 s net130 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X36 VDD net130 Q VDD LPPFET W=0.76U L=0.12U M=1 
X37 Q net130 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X38 VDD net145 c VDD LPPFET W=0.76U L=0.12U M=1 
X39 c net145 VSS VSS LPNFET W=0.28U L=0.12U M=1 
X4 m pm hnet33 VSS LPNFET W=0.5U L=0.12U M=1 
X40 VDD CK net145 VDD LPPFET W=0.28U L=0.12U M=1 
X41 net145 CK VSS VSS LPNFET W=0.28U L=0.12U M=1 
X5 VDD c hnet37 VDD LPPFET W=0.46U L=0.12U M=1 
X6 hnet37 nmin pm VDD LPPFET W=0.46U L=0.12U M=1 
X7 VDD nmset hnet41 VDD LPPFET W=0.28U L=0.12U M=1 
X8 hnet41 RN m VDD LPPFET W=0.28U L=0.12U M=1 
X9 VDD RN hnet45 VDD LPPFET W=0.26U L=0.12U M=1 
.ENDS DFFSRHQX1TS 

**** 
*.SUBCKT DFFSRHQX2TS Q CK D RN SN 
.SUBCKT DFFSRHQX2TS Q CK D RN SN VSS VDD
X0 hnet29 SN VSS VSS LPNFET W=0.84U L=0.12U M=1 
X1 hnet24 cn hnet29 VSS LPNFET W=0.84U L=0.12U M=1 
X10 hnet45 nmset net130 VDD LPPFET W=0.46U L=0.12U M=1 
X11 net90 CK VDD VDD LPPFET W=0.86U L=0.12U M=1 
X12 cn c net90 VDD LPPFET W=0.64U L=0.12U M=1 
X13 pm SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X14 m pm VDD VDD LPPFET W=1.04U L=0.12U M=1 
X15 net100 nmset net99 VDD LPPFET W=0.28U L=0.12U M=1 
X16 net130 c net100 VDD LPPFET W=0.28U L=0.12U M=1 
X17 net99 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X18 net130 cn m VDD LPPFET W=1.14U L=0.12U M=1 
X19 cn CK VSS VSS LPNFET W=0.24U L=0.12U M=1 
X2 pm nmin hnet24 VSS LPNFET W=0.84U L=0.12U M=1 
X20 net115 RN net114 VSS LPNFET W=0.2U L=0.12U M=1 
X21 net130 cn net115 VSS LPNFET W=0.2U L=0.12U M=1 
X22 net114 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X23 net130 nmset VSS VSS LPNFET W=0.2U L=0.12U M=1 
X24 m nmset VSS VSS LPNFET W=0.2U L=0.12U M=1 
X25 net130 c m VSS LPNFET W=0.82U L=0.12U M=1 
X26 hnet47 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X27 pm c hnet47 VSS LPNFET W=0.2U L=0.12U M=1 
X28 hnet49 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X29 VDD m hnet49 VDD LPPFET W=0.28U L=0.12U M=1 
X3 hnet33 RN VSS VSS LPNFET W=0.86U L=0.12U M=1 
X30 VDD SN nmset VDD LPPFET W=0.28U L=0.12U M=1 
X31 nmset SN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X32 VDD D nmin VDD LPPFET W=0.34U L=0.12U M=1 
X33 nmin D VSS VSS LPNFET W=0.24U L=0.12U M=1 
X34 VDD net130 s VDD LPPFET W=0.28U L=0.12U M=1 
X35 s net130 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X36 VDD net130 Q VDD LPPFET W=1.48U L=0.12U M=1 
X37 Q net130 VSS VSS LPNFET W=0.84U L=0.12U M=1 
X38 VDD net145 c VDD LPPFET W=1.12U L=0.12U M=1 
X39 c net145 VSS VSS LPNFET W=0.4U L=0.12U M=1 
X4 m pm hnet33 VSS LPNFET W=0.86U L=0.12U M=1 
X40 VDD CK net145 VDD LPPFET W=0.3U L=0.12U M=1 
X41 net145 CK VSS VSS LPNFET W=0.3U L=0.12U M=1 
X5 VDD c hnet37 VDD LPPFET W=0.8U L=0.12U M=1 
X6 hnet37 nmin pm VDD LPPFET W=0.8U L=0.12U M=1 
X7 VDD nmset hnet41 VDD LPPFET W=0.28U L=0.12U M=1 
X8 hnet41 RN m VDD LPPFET W=0.28U L=0.12U M=1 
X9 VDD RN hnet45 VDD LPPFET W=0.46U L=0.12U M=1 
.ENDS DFFSRHQX2TS 

**** 
*.SUBCKT DFFSRHQX4TS Q CK D RN SN 
.SUBCKT DFFSRHQX4TS Q CK D RN SN VSS VDD
X0 hnet29 RN VSS VSS LPNFET W=0.54U L=0.12U M=1 
X1 m pm hnet29 VSS LPNFET W=0.54U L=0.12U M=1 
X10 pm nmin hnet35 VSS LPNFET W=1.22U L=0.12U M=1 
X11 VDD nmset hnet44 VDD LPPFET W=0.52U L=0.12U M=1 
X12 hnet44 RN m VDD LPPFET W=0.52U L=0.12U M=1 
X13 VDD RN hnet48 VDD LPPFET W=0.84U L=0.12U M=1 
X14 hnet48 nmset net137 VDD LPPFET W=0.84U L=0.12U M=1 
X15 cn c net88 VDD LPPFET W=0.56U L=0.12U M=1 
X16 net88 CK VDD VDD LPPFET W=0.74U L=0.12U M=1 
X17 net97 CK VDD VDD LPPFET W=0.74U L=0.12U M=1 
X18 cn c net97 VDD LPPFET W=0.56U L=0.12U M=1 
X19 pm SN VDD VDD LPPFET W=0.36U L=0.12U M=1 
X2 hnet25 RN VSS VSS LPNFET W=0.54U L=0.12U M=1 
X20 m pm VDD VDD LPPFET W=2.08U L=0.12U M=1 
X21 net109 nmset net113 VDD LPPFET W=0.28U L=0.12U M=1 
X22 net137 c net109 VDD LPPFET W=0.28U L=0.12U M=1 
X23 net113 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X24 net137 cn m VDD LPPFET W=1.3U L=0.12U M=1 
X25 cn CK VSS VSS LPNFET W=0.42U L=0.12U M=1 
X26 net122 RN net121 VSS LPNFET W=0.2U L=0.12U M=1 
X27 net137 cn net122 VSS LPNFET W=0.2U L=0.12U M=1 
X28 net121 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X29 net137 nmset VSS VSS LPNFET W=0.38U L=0.12U M=1 
X3 m pm hnet25 VSS LPNFET W=0.54U L=0.12U M=1 
X30 m nmset VSS VSS LPNFET W=0.38U L=0.12U M=1 
X31 net137 c m VSS LPNFET W=0.92U L=0.12U M=1 
X32 hnet50 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X33 pm c hnet50 VSS LPNFET W=0.2U L=0.12U M=1 
X34 hnet52 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X35 VDD m hnet52 VDD LPPFET W=0.28U L=0.12U M=1 
X36 VDD SN nmset VDD LPPFET W=0.34U L=0.12U M=1 
X37 nmset SN VSS VSS LPNFET W=0.24U L=0.12U M=1 
X38 VDD D nmin VDD LPPFET W=0.62U L=0.12U M=1 
X39 nmin D VSS VSS LPNFET W=0.44U L=0.12U M=1 
X4 VDD c hnet34 VDD LPPFET W=0.6U L=0.12U M=1 
X40 VDD net137 s VDD LPPFET W=0.28U L=0.12U M=1 
X41 s net137 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X42 VDD net137 Q VDD LPPFET W=2.6U L=0.12U M=1 
X43 Q net137 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X44 VDD net152 c VDD LPPFET W=1.84U L=0.12U M=1 
X45 c net152 VSS VSS LPNFET W=0.66U L=0.12U M=1 
X46 VDD CK net152 VDD LPPFET W=0.5U L=0.12U M=1 
X47 net152 CK VSS VSS LPNFET W=0.5U L=0.12U M=1 
X5 hnet34 nmin pm VDD LPPFET W=0.6U L=0.12U M=1 
X6 VDD c hnet31 VDD LPPFET W=0.6U L=0.12U M=1 
X7 hnet31 nmin pm VDD LPPFET W=0.6U L=0.12U M=1 
X8 hnet40 SN VSS VSS LPNFET W=1.22U L=0.12U M=1 
X9 hnet35 cn hnet40 VSS LPNFET W=1.22U L=0.12U M=1 
.ENDS DFFSRHQX4TS 

**** 
*.SUBCKT DFFSRHQX8TS Q CK D RN SN 
.SUBCKT DFFSRHQX8TS Q CK D RN SN VSS VDD
X0 hnet29 RN VSS VSS LPNFET W=0.54U L=0.12U M=1 
X1 m pm hnet29 VSS LPNFET W=0.54U L=0.12U M=1 
X10 pm nmin hnet35 VSS LPNFET W=1.22U L=0.12U M=1 
X11 VDD nmset hnet44 VDD LPPFET W=0.52U L=0.12U M=1 
X12 hnet44 RN m VDD LPPFET W=0.52U L=0.12U M=1 
X13 VDD RN hnet48 VDD LPPFET W=0.84U L=0.12U M=1 
X14 hnet48 nmset net137 VDD LPPFET W=0.84U L=0.12U M=1 
X15 cn c net88 VDD LPPFET W=0.56U L=0.12U M=1 
X16 net88 CK VDD VDD LPPFET W=0.74U L=0.12U M=1 
X17 net97 CK VDD VDD LPPFET W=0.74U L=0.12U M=1 
X18 cn c net97 VDD LPPFET W=0.56U L=0.12U M=1 
X19 pm SN VDD VDD LPPFET W=0.36U L=0.12U M=1 
X2 hnet25 RN VSS VSS LPNFET W=0.54U L=0.12U M=1 
X20 m pm VDD VDD LPPFET W=2.08U L=0.12U M=1 
X21 net109 nmset net113 VDD LPPFET W=0.28U L=0.12U M=1 
X22 net137 c net109 VDD LPPFET W=0.28U L=0.12U M=1 
X23 net113 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X24 net137 cn m VDD LPPFET W=1.3U L=0.12U M=1 
X25 cn CK VSS VSS LPNFET W=0.42U L=0.12U M=1 
X26 net122 RN net121 VSS LPNFET W=0.2U L=0.12U M=1 
X27 net137 cn net122 VSS LPNFET W=0.2U L=0.12U M=1 
X28 net121 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X29 net137 nmset VSS VSS LPNFET W=0.38U L=0.12U M=1 
X3 m pm hnet25 VSS LPNFET W=0.54U L=0.12U M=1 
X30 m nmset VSS VSS LPNFET W=0.38U L=0.12U M=1 
X31 net137 c m VSS LPNFET W=0.92U L=0.12U M=1 
X32 hnet50 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X33 pm c hnet50 VSS LPNFET W=0.2U L=0.12U M=1 
X34 hnet52 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X35 VDD m hnet52 VDD LPPFET W=0.28U L=0.12U M=1 
X36 VDD SN nmset VDD LPPFET W=0.34U L=0.12U M=1 
X37 nmset SN VSS VSS LPNFET W=0.24U L=0.12U M=1 
X38 VDD D nmin VDD LPPFET W=0.62U L=0.12U M=1 
X39 nmin D VSS VSS LPNFET W=0.44U L=0.12U M=1 
X4 VDD c hnet34 VDD LPPFET W=0.6U L=0.12U M=1 
X40 VDD net137 s VDD LPPFET W=0.28U L=0.12U M=1 
X41 s net137 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X42 VDD net137 Q VDD LPPFET W=5.2U L=0.12U M=1 
X43 Q net137 VSS VSS LPNFET W=3.68U L=0.12U M=1 
X44 VDD net152 c VDD LPPFET W=1.84U L=0.12U M=1 
X45 c net152 VSS VSS LPNFET W=0.66U L=0.12U M=1 
X46 VDD CK net152 VDD LPPFET W=0.5U L=0.12U M=1 
X47 net152 CK VSS VSS LPNFET W=0.5U L=0.12U M=1 
X5 hnet34 nmin pm VDD LPPFET W=0.6U L=0.12U M=1 
X6 VDD c hnet31 VDD LPPFET W=0.6U L=0.12U M=1 
X7 hnet31 nmin pm VDD LPPFET W=0.6U L=0.12U M=1 
X8 hnet40 SN VSS VSS LPNFET W=1.22U L=0.12U M=1 
X9 hnet35 cn hnet40 VSS LPNFET W=1.22U L=0.12U M=1 
.ENDS DFFSRHQX8TS 

**** 
*.SUBCKT DFFSRX1TS Q QN CK D RN SN 
.SUBCKT DFFSRX1TS Q QN CK D RN SN VSS VDD
X0 m SN VDD VDD LPPFET W=0.26U L=0.12U M=1 
X1 m pm net64 VDD LPPFET W=0.42U L=0.12U M=1 
X10 net92 s net95 VSS LPNFET W=0.2U L=0.12U M=1 
X11 net95 SN VSS VSS LPNFET W=0.4U L=0.12U M=1 
X12 net101 cn net92 VSS LPNFET W=0.2U L=0.12U M=1 
X13 net101 c m VSS LPNFET W=0.2U L=0.12U M=1 
X14 hnet24 D VSS VSS LPNFET W=0.2U L=0.12U M=1 
X15 pm cn hnet24 VSS LPNFET W=0.2U L=0.12U M=1 
X16 hnet26 c pm VDD LPPFET W=0.28U L=0.12U M=1 
X17 VDD D hnet26 VDD LPPFET W=0.28U L=0.12U M=1 
X18 hnet30 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X19 pm c hnet30 VSS LPNFET W=0.2U L=0.12U M=1 
X2 net64 net114 VDD VDD LPPFET W=0.56U L=0.12U M=1 
X20 hnet32 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X21 VDD m hnet32 VDD LPPFET W=0.28U L=0.12U M=1 
X22 VDD s net110 VDD LPPFET W=0.28U L=0.12U M=1 
X23 net110 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X24 VDD s Q VDD LPPFET W=0.64U L=0.12U M=1 
X25 Q s VSS VSS LPNFET W=0.46U L=0.12U M=1 
X26 VDD RN net114 VDD LPPFET W=0.28U L=0.12U M=1 
X27 net114 RN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X28 VDD net101 s VDD LPPFET W=0.28U L=0.12U M=1 
X29 s net101 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 net101 SN VDD VDD LPPFET W=0.26U L=0.12U M=1 
X30 VDD net110 QN VDD LPPFET W=0.64U L=0.12U M=1 
X31 QN net110 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X32 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X33 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X34 VDD CK cn VDD LPPFET W=0.42U L=0.12U M=1 
X35 cn CK VSS VSS LPNFET W=0.3U L=0.12U M=1 
X4 net74 s net64 VDD LPPFET W=0.28U L=0.12U M=1 
X5 net101 c net74 VDD LPPFET W=0.28U L=0.12U M=1 
X6 net101 cn m VDD LPPFET W=0.28U L=0.12U M=1 
X7 m net114 net95 VSS LPNFET W=0.2U L=0.12U M=1 
X8 m pm net95 VSS LPNFET W=0.3U L=0.12U M=1 
X9 net101 net114 net95 VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS DFFSRX1TS 

**** 
*.SUBCKT DFFSRX2TS Q QN CK D RN SN 
.SUBCKT DFFSRX2TS Q QN CK D RN SN VSS VDD
X0 m SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X1 m pm net62 VDD LPPFET W=0.42U L=0.12U M=1 
X10 net90 s net93 VSS LPNFET W=0.2U L=0.12U M=1 
X11 net93 SN VSS VSS LPNFET W=0.4U L=0.12U M=1 
X12 net99 cn net90 VSS LPNFET W=0.2U L=0.12U M=1 
X13 net99 c m VSS LPNFET W=0.2U L=0.12U M=1 
X14 hnet24 D VSS VSS LPNFET W=0.2U L=0.12U M=1 
X15 pm cn hnet24 VSS LPNFET W=0.2U L=0.12U M=1 
X16 hnet26 c pm VDD LPPFET W=0.28U L=0.12U M=1 
X17 VDD D hnet26 VDD LPPFET W=0.28U L=0.12U M=1 
X18 hnet30 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X19 pm c hnet30 VSS LPNFET W=0.2U L=0.12U M=1 
X2 net62 net112 VDD VDD LPPFET W=0.56U L=0.12U M=1 
X20 hnet32 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X21 VDD m hnet32 VDD LPPFET W=0.28U L=0.12U M=1 
X22 VDD s net108 VDD LPPFET W=0.3U L=0.12U M=1 
X23 net108 s VSS VSS LPNFET W=0.22U L=0.12U M=1 
X24 VDD s Q VDD LPPFET W=1.28U L=0.12U M=1 
X25 Q s VSS VSS LPNFET W=0.92U L=0.12U M=1 
X26 VDD RN net112 VDD LPPFET W=0.28U L=0.12U M=1 
X27 net112 RN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X28 VDD net99 s VDD LPPFET W=0.36U L=0.12U M=1 
X29 s net99 VSS VSS LPNFET W=0.28U L=0.12U M=1 
X3 net99 SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X30 VDD net108 QN VDD LPPFET W=1.28U L=0.12U M=1 
X31 QN net108 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X32 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X33 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X34 VDD CK cn VDD LPPFET W=0.42U L=0.12U M=1 
X35 cn CK VSS VSS LPNFET W=0.3U L=0.12U M=1 
X4 net72 s net62 VDD LPPFET W=0.28U L=0.12U M=1 
X5 net99 c net72 VDD LPPFET W=0.28U L=0.12U M=1 
X6 net99 cn m VDD LPPFET W=0.28U L=0.12U M=1 
X7 m net112 net93 VSS LPNFET W=0.2U L=0.12U M=1 
X8 m pm net93 VSS LPNFET W=0.3U L=0.12U M=1 
X9 net99 net112 net93 VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS DFFSRX2TS 

**** 
*.SUBCKT DFFSRX4TS Q QN CK D RN SN 
.SUBCKT DFFSRX4TS Q QN CK D RN SN VSS VDD
X0 m SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X1 m pm net62 VDD LPPFET W=0.46U L=0.12U M=1 
X10 net90 s net93 VSS LPNFET W=0.2U L=0.12U M=1 
X11 net93 SN VSS VSS LPNFET W=0.46U L=0.12U M=1 
X12 net99 cn net90 VSS LPNFET W=0.2U L=0.12U M=1 
X13 net99 c m VSS LPNFET W=0.22U L=0.12U M=1 
X14 hnet24 D VSS VSS LPNFET W=0.2U L=0.12U M=1 
X15 pm cn hnet24 VSS LPNFET W=0.2U L=0.12U M=1 
X16 hnet26 c pm VDD LPPFET W=0.28U L=0.12U M=1 
X17 VDD D hnet26 VDD LPPFET W=0.28U L=0.12U M=1 
X18 hnet30 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X19 pm c hnet30 VSS LPNFET W=0.2U L=0.12U M=1 
X2 net62 net112 VDD VDD LPPFET W=0.62U L=0.12U M=1 
X20 hnet32 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X21 VDD m hnet32 VDD LPPFET W=0.28U L=0.12U M=1 
X22 VDD s net108 VDD LPPFET W=0.62U L=0.12U M=1 
X23 net108 s VSS VSS LPNFET W=0.4U L=0.12U M=1 
X24 VDD s Q VDD LPPFET W=2.4U L=0.12U M=1 
X25 Q s VSS VSS LPNFET W=1.84U L=0.12U M=1 
X26 VDD RN net112 VDD LPPFET W=0.28U L=0.12U M=1 
X27 net112 RN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X28 VDD net99 s VDD LPPFET W=0.66U L=0.12U M=1 
X29 s net99 VSS VSS LPNFET W=0.44U L=0.12U M=1 
X3 net99 SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X30 VDD net108 QN VDD LPPFET W=2.4U L=0.12U M=1 
X31 QN net108 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X32 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X33 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X34 VDD CK cn VDD LPPFET W=0.44U L=0.12U M=1 
X35 cn CK VSS VSS LPNFET W=0.32U L=0.12U M=1 
X4 net72 s net62 VDD LPPFET W=0.28U L=0.12U M=1 
X5 net99 c net72 VDD LPPFET W=0.28U L=0.12U M=1 
X6 net99 cn m VDD LPPFET W=0.3U L=0.12U M=1 
X7 m net112 net93 VSS LPNFET W=0.2U L=0.12U M=1 
X8 m pm net93 VSS LPNFET W=0.34U L=0.12U M=1 
X9 net99 net112 net93 VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS DFFSRX4TS 

**** 
*.SUBCKT DFFSRXLTS Q QN CK D RN SN 
.SUBCKT DFFSRXLTS Q QN CK D RN SN VSS VDD
X0 m SN VDD VDD LPPFET W=0.26U L=0.12U M=1 
X1 m pm net62 VDD LPPFET W=0.42U L=0.12U M=1 
X10 net90 s net93 VSS LPNFET W=0.2U L=0.12U M=1 
X11 net93 SN VSS VSS LPNFET W=0.4U L=0.12U M=1 
X12 net99 cn net90 VSS LPNFET W=0.2U L=0.12U M=1 
X13 net99 c m VSS LPNFET W=0.2U L=0.12U M=1 
X14 hnet24 D VSS VSS LPNFET W=0.2U L=0.12U M=1 
X15 pm cn hnet24 VSS LPNFET W=0.2U L=0.12U M=1 
X16 hnet26 c pm VDD LPPFET W=0.28U L=0.12U M=1 
X17 VDD D hnet26 VDD LPPFET W=0.28U L=0.12U M=1 
X18 hnet30 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X19 pm c hnet30 VSS LPNFET W=0.2U L=0.12U M=1 
X2 net62 net112 VDD VDD LPPFET W=0.56U L=0.12U M=1 
X20 hnet32 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X21 VDD m hnet32 VDD LPPFET W=0.28U L=0.12U M=1 
X22 VDD s net108 VDD LPPFET W=0.28U L=0.12U M=1 
X23 net108 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X24 VDD s Q VDD LPPFET W=0.34U L=0.12U M=1 
X25 Q s VSS VSS LPNFET W=0.24U L=0.12U M=1 
X26 VDD RN net112 VDD LPPFET W=0.28U L=0.12U M=1 
X27 net112 RN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X28 VDD net99 s VDD LPPFET W=0.28U L=0.12U M=1 
X29 s net99 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 net99 SN VDD VDD LPPFET W=0.26U L=0.12U M=1 
X30 VDD net108 QN VDD LPPFET W=0.34U L=0.12U M=1 
X31 QN net108 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X32 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X33 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X34 VDD CK cn VDD LPPFET W=0.42U L=0.12U M=1 
X35 cn CK VSS VSS LPNFET W=0.3U L=0.12U M=1 
X4 net72 s net62 VDD LPPFET W=0.28U L=0.12U M=1 
X5 net99 c net72 VDD LPPFET W=0.28U L=0.12U M=1 
X6 net99 cn m VDD LPPFET W=0.28U L=0.12U M=1 
X7 m net112 net93 VSS LPNFET W=0.2U L=0.12U M=1 
X8 m pm net93 VSS LPNFET W=0.3U L=0.12U M=1 
X9 net99 net112 net93 VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS DFFSRXLTS 

**** 
*.SUBCKT DFFSX1TS Q QN CK D SN 
.SUBCKT DFFSX1TS Q QN CK D SN VSS VDD
X0 net52 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X1 m SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X10 net82 c m VSS LPNFET W=0.2U L=0.12U M=1 
X11 hnet21 D VSS VSS LPNFET W=0.2U L=0.12U M=1 
X12 pm cn hnet21 VSS LPNFET W=0.2U L=0.12U M=1 
X13 hnet23 c pm VDD LPPFET W=0.28U L=0.12U M=1 
X14 VDD D hnet23 VDD LPPFET W=0.28U L=0.12U M=1 
X15 hnet27 m VSS VSS LPNFET W=0.22U L=0.12U M=1 
X16 pm c hnet27 VSS LPNFET W=0.22U L=0.12U M=1 
X17 hnet29 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X18 VDD m hnet29 VDD LPPFET W=0.28U L=0.12U M=1 
X19 VDD s net91 VDD LPPFET W=0.28U L=0.12U M=1 
X2 m pm VDD VDD LPPFET W=0.28U L=0.12U M=1 
X20 net91 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X21 VDD s Q VDD LPPFET W=0.64U L=0.12U M=1 
X22 Q s VSS VSS LPNFET W=0.46U L=0.12U M=1 
X23 VDD net82 s VDD LPPFET W=0.28U L=0.12U M=1 
X24 s net82 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X25 VDD net91 QN VDD LPPFET W=0.64U L=0.12U M=1 
X26 QN net91 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X27 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X28 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X29 VDD CK cn VDD LPPFET W=0.42U L=0.12U M=1 
X3 net82 SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X30 cn CK VSS VSS LPNFET W=0.3U L=0.12U M=1 
X4 net82 c net52 VDD LPPFET W=0.28U L=0.12U M=1 
X5 net82 cn m VDD LPPFET W=0.28U L=0.12U M=1 
X6 m pm net76 VSS LPNFET W=0.3U L=0.12U M=1 
X7 net73 s net76 VSS LPNFET W=0.2U L=0.12U M=1 
X8 net76 SN VSS VSS LPNFET W=0.4U L=0.12U M=1 
X9 net82 cn net73 VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS DFFSX1TS 

**** 
*.SUBCKT DFFSX2TS Q QN CK D SN 
.SUBCKT DFFSX2TS Q QN CK D SN VSS VDD
X0 net52 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X1 m SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X10 net82 c m VSS LPNFET W=0.2U L=0.12U M=1 
X11 hnet21 D VSS VSS LPNFET W=0.2U L=0.12U M=1 
X12 pm cn hnet21 VSS LPNFET W=0.2U L=0.12U M=1 
X13 hnet23 c pm VDD LPPFET W=0.28U L=0.12U M=1 
X14 VDD D hnet23 VDD LPPFET W=0.28U L=0.12U M=1 
X15 hnet27 m VSS VSS LPNFET W=0.22U L=0.12U M=1 
X16 pm c hnet27 VSS LPNFET W=0.22U L=0.12U M=1 
X17 hnet29 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X18 VDD m hnet29 VDD LPPFET W=0.28U L=0.12U M=1 
X19 VDD s net91 VDD LPPFET W=0.3U L=0.12U M=1 
X2 m pm VDD VDD LPPFET W=0.28U L=0.12U M=1 
X20 net91 s VSS VSS LPNFET W=0.22U L=0.12U M=1 
X21 VDD s Q VDD LPPFET W=1.28U L=0.12U M=1 
X22 Q s VSS VSS LPNFET W=0.92U L=0.12U M=1 
X23 VDD net82 s VDD LPPFET W=0.34U L=0.12U M=1 
X24 s net82 VSS VSS LPNFET W=0.26U L=0.12U M=1 
X25 VDD net91 QN VDD LPPFET W=1.28U L=0.12U M=1 
X26 QN net91 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X27 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X28 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X29 VDD CK cn VDD LPPFET W=0.42U L=0.12U M=1 
X3 net82 SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X30 cn CK VSS VSS LPNFET W=0.3U L=0.12U M=1 
X4 net82 c net52 VDD LPPFET W=0.28U L=0.12U M=1 
X5 net82 cn m VDD LPPFET W=0.28U L=0.12U M=1 
X6 m pm net76 VSS LPNFET W=0.3U L=0.12U M=1 
X7 net73 s net76 VSS LPNFET W=0.2U L=0.12U M=1 
X8 net76 SN VSS VSS LPNFET W=0.4U L=0.12U M=1 
X9 net82 cn net73 VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS DFFSX2TS 

**** 
*.SUBCKT DFFSX4TS Q QN CK D SN 
.SUBCKT DFFSX4TS Q QN CK D SN VSS VDD
X0 net52 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X1 m SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X10 net82 c m VSS LPNFET W=0.24U L=0.12U M=1 
X11 hnet21 D VSS VSS LPNFET W=0.2U L=0.12U M=1 
X12 pm cn hnet21 VSS LPNFET W=0.2U L=0.12U M=1 
X13 hnet23 c pm VDD LPPFET W=0.28U L=0.12U M=1 
X14 VDD D hnet23 VDD LPPFET W=0.28U L=0.12U M=1 
X15 hnet27 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X16 pm c hnet27 VSS LPNFET W=0.2U L=0.12U M=1 
X17 hnet29 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X18 VDD m hnet29 VDD LPPFET W=0.28U L=0.12U M=1 
X19 VDD s net91 VDD LPPFET W=0.62U L=0.12U M=1 
X2 m pm VDD VDD LPPFET W=0.34U L=0.12U M=1 
X20 net91 s VSS VSS LPNFET W=0.44U L=0.12U M=1 
X21 VDD s Q VDD LPPFET W=2.56U L=0.12U M=1 
X22 Q s VSS VSS LPNFET W=1.84U L=0.12U M=1 
X23 VDD net82 s VDD LPPFET W=0.7U L=0.12U M=1 
X24 s net82 VSS VSS LPNFET W=0.5U L=0.12U M=1 
X25 VDD net91 QN VDD LPPFET W=2.56U L=0.12U M=1 
X26 QN net91 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X27 VDD cn c VDD LPPFET W=0.3U L=0.12U M=1 
X28 c cn VSS VSS LPNFET W=0.22U L=0.12U M=1 
X29 VDD CK cn VDD LPPFET W=0.44U L=0.12U M=1 
X3 net82 SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X30 cn CK VSS VSS LPNFET W=0.32U L=0.12U M=1 
X4 net82 c net52 VDD LPPFET W=0.28U L=0.12U M=1 
X5 net82 cn m VDD LPPFET W=0.34U L=0.12U M=1 
X6 m pm net76 VSS LPNFET W=0.36U L=0.12U M=1 
X7 net73 s net76 VSS LPNFET W=0.2U L=0.12U M=1 
X8 net76 SN VSS VSS LPNFET W=0.48U L=0.12U M=1 
X9 net82 cn net73 VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS DFFSX4TS 

**** 
*.SUBCKT DFFSXLTS Q QN CK D SN 
.SUBCKT DFFSXLTS Q QN CK D SN VSS VDD
X0 net52 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X1 m SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X10 net82 c m VSS LPNFET W=0.2U L=0.12U M=1 
X11 hnet21 D VSS VSS LPNFET W=0.2U L=0.12U M=1 
X12 pm cn hnet21 VSS LPNFET W=0.2U L=0.12U M=1 
X13 hnet23 c pm VDD LPPFET W=0.28U L=0.12U M=1 
X14 VDD D hnet23 VDD LPPFET W=0.28U L=0.12U M=1 
X15 hnet27 m VSS VSS LPNFET W=0.22U L=0.12U M=1 
X16 pm c hnet27 VSS LPNFET W=0.22U L=0.12U M=1 
X17 hnet29 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X18 VDD m hnet29 VDD LPPFET W=0.28U L=0.12U M=1 
X19 VDD s net91 VDD LPPFET W=0.28U L=0.12U M=1 
X2 m pm VDD VDD LPPFET W=0.28U L=0.12U M=1 
X20 net91 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X21 VDD s Q VDD LPPFET W=0.34U L=0.12U M=1 
X22 Q s VSS VSS LPNFET W=0.24U L=0.12U M=1 
X23 VDD net82 s VDD LPPFET W=0.28U L=0.12U M=1 
X24 s net82 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X25 VDD net91 QN VDD LPPFET W=0.34U L=0.12U M=1 
X26 QN net91 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X27 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X28 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X29 VDD CK cn VDD LPPFET W=0.42U L=0.12U M=1 
X3 net82 SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X30 cn CK VSS VSS LPNFET W=0.3U L=0.12U M=1 
X4 net82 c net52 VDD LPPFET W=0.28U L=0.12U M=1 
X5 net82 cn m VDD LPPFET W=0.28U L=0.12U M=1 
X6 m pm net76 VSS LPNFET W=0.3U L=0.12U M=1 
X7 net73 s net76 VSS LPNFET W=0.2U L=0.12U M=1 
X8 net76 SN VSS VSS LPNFET W=0.4U L=0.12U M=1 
X9 net82 cn net73 VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS DFFSXLTS 

**** 
*.SUBCKT DFFTRX1TS Q QN CK D RN 
.SUBCKT DFFTRX1TS Q QN CK D RN VSS VDD
X0 VDD m hnet23 VDD LPPFET W=0.28U L=0.12U M=1 
X1 hnet23 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X10 net83 c net67 VDD LPPFET W=0.28U L=0.12U M=1 
X11 net67 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X12 net83 cn m VDD LPPFET W=0.28U L=0.12U M=1 
X13 net83 cn net80 VSS LPNFET W=0.2U L=0.12U M=1 
X14 net80 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X15 net83 c m VSS LPNFET W=0.2U L=0.12U M=1 
X16 VDD s net84 VDD LPPFET W=0.28U L=0.12U M=1 
X17 net84 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X18 VDD net83 s VDD LPPFET W=0.28U L=0.12U M=1 
X19 s net83 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 hnet27 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X20 VDD pm m VDD LPPFET W=0.28U L=0.12U M=1 
X21 m pm VSS VSS LPNFET W=0.2U L=0.12U M=1 
X22 VDD s Q VDD LPPFET W=0.64U L=0.12U M=1 
X23 Q s VSS VSS LPNFET W=0.46U L=0.12U M=1 
X24 VDD net84 QN VDD LPPFET W=0.64U L=0.12U M=1 
X25 QN net84 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X26 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X27 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X28 VDD CK cn VDD LPPFET W=0.42U L=0.12U M=1 
X29 cn CK VSS VSS LPNFET W=0.3U L=0.12U M=1 
X3 pm c hnet27 VSS LPNFET W=0.2U L=0.12U M=1 
X4 hnet33 RN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X5 hnet28 D hnet33 VSS LPNFET W=0.2U L=0.12U M=1 
X6 pm cn hnet28 VSS LPNFET W=0.2U L=0.12U M=1 
X7 net64 RN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X8 net64 D VDD VDD LPPFET W=0.28U L=0.12U M=1 
X9 pm c net64 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS DFFTRX1TS 

****.SUBCKT DFFTRX2TS Q QN CK D RN 
*.SUBCKT DFFTRX2TS CK D Q QN RN 
.SUBCKT DFFTRX2TS CK D Q QN RN VSS VDD
X0 VDD m hnet23 VDD LPPFET W=0.28U L=0.12U M=1 
X1 hnet23 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X10 net83 c net67 VDD LPPFET W=0.28U L=0.12U M=1 
X11 net67 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X12 net83 cn m VDD LPPFET W=0.28U L=0.12U M=1 
X13 net83 cn net80 VSS LPNFET W=0.2U L=0.12U M=1 
X14 net80 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X15 net83 c m VSS LPNFET W=0.2U L=0.12U M=1 
X16 VDD s net84 VDD LPPFET W=0.3U L=0.12U M=1 
X17 net84 s VSS VSS LPNFET W=0.22U L=0.12U M=1 
X18 VDD net83 s VDD LPPFET W=0.36U L=0.12U M=1 
X19 s net83 VSS VSS LPNFET W=0.26U L=0.12U M=1 
X2 hnet27 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X20 VDD pm m VDD LPPFET W=0.28U L=0.12U M=1 
X21 m pm VSS VSS LPNFET W=0.2U L=0.12U M=1 
X22 VDD s Q VDD LPPFET W=1.28U L=0.12U M=1 
X23 Q s VSS VSS LPNFET W=0.92U L=0.12U M=1 
X24 VDD net84 QN VDD LPPFET W=1.28U L=0.12U M=1 
X25 QN net84 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X26 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X27 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X28 VDD CK cn VDD LPPFET W=0.42U L=0.12U M=1 
X29 cn CK VSS VSS LPNFET W=0.3U L=0.12U M=1 
X3 pm c hnet27 VSS LPNFET W=0.2U L=0.12U M=1 
X4 hnet33 RN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X5 hnet28 D hnet33 VSS LPNFET W=0.2U L=0.12U M=1 
X6 pm cn hnet28 VSS LPNFET W=0.2U L=0.12U M=1 
X7 net64 RN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X8 net64 D VDD VDD LPPFET W=0.28U L=0.12U M=1 
X9 pm c net64 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS DFFTRX2TS 

**** 
*.SUBCKT DFFTRX4TS Q QN CK D RN 
.SUBCKT DFFTRX4TS Q QN CK D RN VSS VDD
X0 VDD m hnet23 VDD LPPFET W=0.28U L=0.12U M=1 
X1 hnet23 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X10 net83 c net67 VDD LPPFET W=0.28U L=0.12U M=1 
X11 net67 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X12 net83 cn m VDD LPPFET W=0.3U L=0.12U M=1 
X13 net83 cn net80 VSS LPNFET W=0.2U L=0.12U M=1 
X14 net80 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X15 net83 c m VSS LPNFET W=0.22U L=0.12U M=1 
X16 VDD s net84 VDD LPPFET W=0.62U L=0.12U M=1 
X17 net84 s VSS VSS LPNFET W=0.4U L=0.12U M=1 
X18 VDD net83 s VDD LPPFET W=0.66U L=0.12U M=1 
X19 s net83 VSS VSS LPNFET W=0.44U L=0.12U M=1 
X2 hnet27 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X20 VDD pm m VDD LPPFET W=0.3U L=0.12U M=1 
X21 m pm VSS VSS LPNFET W=0.22U L=0.12U M=1 
X22 VDD s Q VDD LPPFET W=2.4U L=0.12U M=1 
X23 Q s VSS VSS LPNFET W=1.84U L=0.12U M=1 
X24 VDD net84 QN VDD LPPFET W=2.4U L=0.12U M=1 
X25 QN net84 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X26 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X27 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X28 VDD CK cn VDD LPPFET W=0.44U L=0.12U M=1 
X29 cn CK VSS VSS LPNFET W=0.32U L=0.12U M=1 
X3 pm c hnet27 VSS LPNFET W=0.2U L=0.12U M=1 
X4 hnet33 RN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X5 hnet28 D hnet33 VSS LPNFET W=0.2U L=0.12U M=1 
X6 pm cn hnet28 VSS LPNFET W=0.2U L=0.12U M=1 
X7 net64 RN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X8 net64 D VDD VDD LPPFET W=0.28U L=0.12U M=1 
X9 pm c net64 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS DFFTRX4TS 

**** 
*.SUBCKT DFFTRXLTS Q QN CK D RN 
.SUBCKT DFFTRXLTS Q QN CK D RN VSS VDD
X0 VDD m hnet23 VDD LPPFET W=0.28U L=0.12U M=1 
X1 hnet23 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X10 net83 c net67 VDD LPPFET W=0.28U L=0.12U M=1 
X11 net67 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X12 net83 cn m VDD LPPFET W=0.28U L=0.12U M=1 
X13 net83 cn net80 VSS LPNFET W=0.2U L=0.12U M=1 
X14 net80 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X15 net83 c m VSS LPNFET W=0.2U L=0.12U M=1 
X16 VDD s net84 VDD LPPFET W=0.28U L=0.12U M=1 
X17 net84 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X18 VDD net83 s VDD LPPFET W=0.28U L=0.12U M=1 
X19 s net83 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 hnet27 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X20 VDD pm m VDD LPPFET W=0.28U L=0.12U M=1 
X21 m pm VSS VSS LPNFET W=0.2U L=0.12U M=1 
X22 VDD s Q VDD LPPFET W=0.34U L=0.12U M=1 
X23 Q s VSS VSS LPNFET W=0.24U L=0.12U M=1 
X24 VDD net84 QN VDD LPPFET W=0.34U L=0.12U M=1 
X25 QN net84 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X26 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X27 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X28 VDD CK cn VDD LPPFET W=0.42U L=0.12U M=1 
X29 cn CK VSS VSS LPNFET W=0.3U L=0.12U M=1 
X3 pm c hnet27 VSS LPNFET W=0.2U L=0.12U M=1 
X4 hnet33 RN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X5 hnet28 D hnet33 VSS LPNFET W=0.2U L=0.12U M=1 
X6 pm cn hnet28 VSS LPNFET W=0.2U L=0.12U M=1 
X7 net64 RN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X8 net64 D VDD VDD LPPFET W=0.28U L=0.12U M=1 
X9 pm c net64 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS DFFTRXLTS 

**** 
*.SUBCKT DFFX1TS Q QN CK D 
.SUBCKT DFFX1TS Q QN CK D VSS VDD
X0 hnet14 m VSS VSS LPNFET W=0.58U L=0.12U M=1 
X1 net43 c hnet14 VSS LPNFET W=0.58U L=0.12U M=1 
X10 hnet32 c net43 VDD LPPFET W=0.28U L=0.12U M=1 
X11 VDD s hnet32 VDD LPPFET W=0.28U L=0.12U M=1 
X12 hnet38 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X13 pm c hnet38 VSS LPNFET W=0.2U L=0.12U M=1 
X14 hnet40 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X15 VDD m hnet40 VDD LPPFET W=0.28U L=0.12U M=1 
X16 VDD net43 s VDD LPPFET W=0.36U L=0.12U M=1 
X17 s net43 VSS VSS LPNFET W=0.26U L=0.12U M=1 
X18 VDD pm m VDD LPPFET W=0.3U L=0.12U M=1 
X19 m pm VSS VSS LPNFET W=0.22U L=0.12U M=1 
X2 hnet16 cn net43 VDD LPPFET W=0.8U L=0.12U M=1 
X20 VDD s QN VDD LPPFET W=0.64U L=0.12U M=1 
X21 QN s VSS VSS LPNFET W=0.46U L=0.12U M=1 
X22 VDD cn c VDD LPPFET W=0.34U L=0.12U M=1 
X23 c cn VSS VSS LPNFET W=0.24U L=0.12U M=1 
X24 VDD CK cn VDD LPPFET W=0.48U L=0.12U M=1 
X25 cn CK VSS VSS LPNFET W=0.34U L=0.12U M=1 
X26 VDD net43 Q VDD LPPFET W=0.64U L=0.12U M=1 
X27 Q net43 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X3 VDD m hnet16 VDD LPPFET W=0.8U L=0.12U M=1 
X4 hnet22 D VSS VSS LPNFET W=0.2U L=0.12U M=1 
X5 pm cn hnet22 VSS LPNFET W=0.2U L=0.12U M=1 
X6 hnet24 c pm VDD LPPFET W=0.28U L=0.12U M=1 
X7 VDD D hnet24 VDD LPPFET W=0.28U L=0.12U M=1 
X8 hnet30 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X9 net43 cn hnet30 VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS DFFX1TS 

**** 
*.SUBCKT DFFX2TS Q QN CK D 
.SUBCKT DFFX2TS Q QN CK D VSS VDD
X0 hnet14 m VSS VSS LPNFET W=0.54U L=0.12U M=1 
X1 hnet15 m VSS VSS LPNFET W=0.54U L=0.12U M=1 
X10 hnet26 c pm VDD LPPFET W=0.38U L=0.12U M=1 
X11 VDD D hnet26 VDD LPPFET W=0.38U L=0.12U M=1 
X12 hnet30 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X13 net43 cn hnet30 VSS LPNFET W=0.2U L=0.12U M=1 
X14 hnet32 c net43 VDD LPPFET W=0.28U L=0.12U M=1 
X15 VDD s hnet32 VDD LPPFET W=0.28U L=0.12U M=1 
X16 hnet36 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X17 pm c hnet36 VSS LPNFET W=0.2U L=0.12U M=1 
X18 hnet38 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X19 VDD m hnet38 VDD LPPFET W=0.28U L=0.12U M=1 
X2 net43 c hnet14 VSS LPNFET W=0.54U L=0.12U M=1 
X20 VDD net43 s VDD LPPFET W=0.62U L=0.12U M=1 
X21 s net43 VSS VSS LPNFET W=0.44U L=0.12U M=1 
X22 VDD pm m VDD LPPFET W=0.5U L=0.12U M=1 
X23 m pm VSS VSS LPNFET W=0.36U L=0.12U M=1 
X24 VDD s QN VDD LPPFET W=1.28U L=0.12U M=1 
X25 QN s VSS VSS LPNFET W=0.92U L=0.12U M=1 
X26 VDD cn c VDD LPPFET W=0.5U L=0.12U M=1 
X27 c cn VSS VSS LPNFET W=0.36U L=0.12U M=1 
X28 VDD CK cn VDD LPPFET W=0.7U L=0.12U M=1 
X29 cn CK VSS VSS LPNFET W=0.5U L=0.12U M=1 
X3 net43 c hnet15 VSS LPNFET W=0.54U L=0.12U M=1 
X30 VDD net43 Q VDD LPPFET W=1.28U L=0.12U M=1 
X31 Q net43 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X4 hnet22 cn net43 VDD LPPFET W=0.76U L=0.12U M=1 
X5 hnet19 cn net43 VDD LPPFET W=0.76U L=0.12U M=1 
X6 VDD m hnet22 VDD LPPFET W=0.76U L=0.12U M=1 
X7 VDD m hnet19 VDD LPPFET W=0.76U L=0.12U M=1 
X8 hnet24 D VSS VSS LPNFET W=0.28U L=0.12U M=1 
X9 pm cn hnet24 VSS LPNFET W=0.28U L=0.12U M=1 
.ENDS DFFX2TS 

**** 
*.SUBCKT DFFX4TS Q QN CK D 
.SUBCKT DFFX4TS Q QN CK D VSS VDD
X0 hnet15 m VSS VSS LPNFET W=0.7U L=0.12U M=1 
X1 hnet17 m VSS VSS LPNFET W=0.7U L=0.12U M=1 
X10 VDD m hnet18 VDD LPPFET W=0.98U L=0.12U M=1 
X11 VDD m hnet14 VDD LPPFET W=0.98U L=0.12U M=1 
X12 hnet26 D VSS VSS LPNFET W=0.52U L=0.12U M=1 
X13 pm cn hnet26 VSS LPNFET W=0.52U L=0.12U M=1 
X14 hnet28 c pm VDD LPPFET W=0.72U L=0.12U M=1 
X15 VDD D hnet28 VDD LPPFET W=0.72U L=0.12U M=1 
X16 hnet32 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X17 net43 cn hnet32 VSS LPNFET W=0.2U L=0.12U M=1 
X18 hnet34 c net43 VDD LPPFET W=0.28U L=0.12U M=1 
X19 VDD s hnet34 VDD LPPFET W=0.28U L=0.12U M=1 
X2 hnet22 m VSS VSS LPNFET W=0.7U L=0.12U M=1 
X20 hnet38 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X21 pm c hnet38 VSS LPNFET W=0.2U L=0.12U M=1 
X22 hnet40 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X23 VDD m hnet40 VDD LPPFET W=0.28U L=0.12U M=1 
X24 VDD net43 s VDD LPPFET W=1.14U L=0.12U M=1 
X25 s net43 VSS VSS LPNFET W=0.82U L=0.12U M=1 
X26 VDD pm m VDD LPPFET W=0.92U L=0.12U M=1 
X27 m pm VSS VSS LPNFET W=0.66U L=0.12U M=1 
X28 VDD s QN VDD LPPFET W=2.56U L=0.12U M=1 
X29 QN s VSS VSS LPNFET W=1.84U L=0.12U M=1 
X3 net43 c hnet15 VSS LPNFET W=0.7U L=0.12U M=1 
X30 VDD cn c VDD LPPFET W=0.84U L=0.12U M=1 
X31 c cn VSS VSS LPNFET W=0.6U L=0.12U M=1 
X32 VDD CK cn VDD LPPFET W=1.12U L=0.12U M=1 
X33 cn CK VSS VSS LPNFET W=0.78U L=0.12U M=1 
X34 VDD net43 Q VDD LPPFET W=2.56U L=0.12U M=1 
X35 Q net43 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X4 net43 c hnet17 VSS LPNFET W=0.7U L=0.12U M=1 
X5 net43 c hnet22 VSS LPNFET W=0.7U L=0.12U M=1 
X6 hnet16 cn net43 VDD LPPFET W=0.98U L=0.12U M=1 
X7 hnet18 cn net43 VDD LPPFET W=0.98U L=0.12U M=1 
X8 hnet14 cn net43 VDD LPPFET W=0.98U L=0.12U M=1 
X9 VDD m hnet16 VDD LPPFET W=0.98U L=0.12U M=1 
.ENDS DFFX4TS 

**** 
*.SUBCKT DFFXLTS Q QN CK D 
.SUBCKT DFFXLTS Q QN CK D VSS VDD
X0 hnet14 m VSS VSS LPNFET W=0.36U L=0.12U M=1 
X1 net43 c hnet14 VSS LPNFET W=0.36U L=0.12U M=1 
X10 hnet32 c net43 VDD LPPFET W=0.28U L=0.12U M=1 
X11 VDD s hnet32 VDD LPPFET W=0.28U L=0.12U M=1 
X12 hnet38 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X13 pm c hnet38 VSS LPNFET W=0.2U L=0.12U M=1 
X14 hnet40 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X15 VDD m hnet40 VDD LPPFET W=0.28U L=0.12U M=1 
X16 VDD net43 s VDD LPPFET W=0.28U L=0.12U M=1 
X17 s net43 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X18 VDD pm m VDD LPPFET W=0.28U L=0.12U M=1 
X19 m pm VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 hnet16 cn net43 VDD LPPFET W=0.5U L=0.12U M=1 
X20 VDD s QN VDD LPPFET W=0.34U L=0.12U M=1 
X21 QN s VSS VSS LPNFET W=0.24U L=0.12U M=1 
X22 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X23 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X24 VDD CK cn VDD LPPFET W=0.38U L=0.12U M=1 
X25 cn CK VSS VSS LPNFET W=0.28U L=0.12U M=1 
X26 VDD net43 Q VDD LPPFET W=0.34U L=0.12U M=1 
X27 Q net43 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X3 VDD m hnet16 VDD LPPFET W=0.5U L=0.12U M=1 
X4 hnet22 D VSS VSS LPNFET W=0.2U L=0.12U M=1 
X5 pm cn hnet22 VSS LPNFET W=0.2U L=0.12U M=1 
X6 hnet24 c pm VDD LPPFET W=0.28U L=0.12U M=1 
X7 VDD D hnet24 VDD LPPFET W=0.28U L=0.12U M=1 
X8 hnet30 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X9 net43 cn hnet30 VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS DFFXLTS 

**** 
*.SUBCKT DLY1X1TS Y A 
.SUBCKT DLY1X1TS Y A VSS VDD
X0 net18 nmin VSS VSS LPNFET W=0.52U L=0.12U M=1 
X1 net21 net18 VSS VSS LPNFET W=0.52U L=0.12U M=1 
X2 net18 nmin VDD VDD LPPFET W=0.8U L=0.12U M=1 
X3 net21 net18 VDD VDD LPPFET W=0.8U L=0.12U M=1 
X4 VDD A nmin VDD LPPFET W=0.8U L=0.12U M=1 
X5 nmin A VSS VSS LPNFET W=0.52U L=0.12U M=1 
X6 VDD net21 Y VDD LPPFET W=0.64U L=0.12U M=1 
X7 Y net21 VSS VSS LPNFET W=0.24U L=0.12U M=1 
.ENDS DLY1X1TS 

**** 
*.SUBCKT DLY1X4TS Y A 
.SUBCKT DLY1X4TS Y A VSS VDD
X0 net18 nmin VSS VSS LPNFET W=0.58U L=0.12U M=1 
X1 net21 net18 VSS VSS LPNFET W=0.58U L=0.12U M=1 
X2 net18 nmin VDD VDD LPPFET W=0.8U L=0.12U M=1 
X3 net21 net18 VDD VDD LPPFET W=0.8U L=0.12U M=1 
X4 VDD A nmin VDD LPPFET W=0.8U L=0.12U M=1 
X5 nmin A VSS VSS LPNFET W=0.58U L=0.12U M=1 
X6 VDD net21 Y VDD LPPFET W=2.54U L=0.12U M=1 
X7 Y net21 VSS VSS LPNFET W=0.92U L=0.12U M=1 
.ENDS DLY1X4TS 

**** 
*.SUBCKT DLY2X1TS Y A 
.SUBCKT DLY2X1TS Y A VSS VDD
X0 net18 nmin VSS VSS LPNFET W=0.52U L=0.24U M=1 
X1 net21 net18 VSS VSS LPNFET W=0.52U L=0.24U M=1 
X2 net18 nmin VDD VDD LPPFET W=0.72U L=0.24U M=1 
X3 net21 net18 VDD VDD LPPFET W=0.72U L=0.24U M=1 
X4 VDD A nmin VDD LPPFET W=0.72U L=0.12U M=1 
X5 nmin A VSS VSS LPNFET W=0.24U L=0.12U M=1 
X6 VDD net21 Y VDD LPPFET W=0.64U L=0.12U M=1 
X7 Y net21 VSS VSS LPNFET W=0.24U L=0.12U M=1 
.ENDS DLY2X1TS 

**** 
*.SUBCKT DLY2X4TS Y A 
.SUBCKT DLY2X4TS Y A VSS VDD
X0 net18 nmin VSS VSS LPNFET W=0.58U L=0.3U M=1 
X1 net21 net18 VSS VSS LPNFET W=0.58U L=0.3U M=1 
X2 net18 nmin VDD VDD LPPFET W=0.8U L=0.3U M=1 
X3 net21 net18 VDD VDD LPPFET W=0.8U L=0.3U M=1 
X4 VDD A nmin VDD LPPFET W=0.8U L=0.12U M=1 
X5 nmin A VSS VSS LPNFET W=0.58U L=0.12U M=1 
X6 VDD net21 Y VDD LPPFET W=2.54U L=0.12U M=1 
X7 Y net21 VSS VSS LPNFET W=0.92U L=0.12U M=1 
.ENDS DLY2X4TS 

**** 
*.SUBCKT DLY3X1TS Y A 
.SUBCKT DLY3X1TS Y A VSS VDD
X0 net18 nmin VSS VSS LPNFET W=0.52U L=0.44U M=1 
X1 net21 net18 VSS VSS LPNFET W=0.52U L=0.44U M=1 
X2 net18 nmin VDD VDD LPPFET W=0.72U L=0.44U M=1 
X3 net21 net18 VDD VDD LPPFET W=0.72U L=0.44U M=1 
X4 VDD A nmin VDD LPPFET W=0.72U L=0.12U M=1 
X5 nmin A VSS VSS LPNFET W=0.52U L=0.12U M=1 
X6 VDD net21 Y VDD LPPFET W=0.64U L=0.12U M=1 
X7 Y net21 VSS VSS LPNFET W=0.24U L=0.12U M=1 
.ENDS DLY3X1TS 

**** 
*.SUBCKT DLY3X4TS Y A 
.SUBCKT DLY3X4TS Y A VSS VDD
X0 net18 nmin VSS VSS LPNFET W=0.58U L=0.48U M=1 
X1 net21 net18 VSS VSS LPNFET W=0.58U L=0.48U M=1 
X2 net18 nmin VDD VDD LPPFET W=0.8U L=0.48U M=1 
X3 net21 net18 VDD VDD LPPFET W=0.8U L=0.48U M=1 
X4 VDD A nmin VDD LPPFET W=0.8U L=0.12U M=1 
X5 nmin A VSS VSS LPNFET W=0.58U L=0.12U M=1 
X6 VDD net21 Y VDD LPPFET W=2.54U L=0.12U M=1 
X7 Y net21 VSS VSS LPNFET W=0.92U L=0.12U M=1 
.ENDS DLY3X4TS 

**** 
*.SUBCKT DLY4X1TS Y A 
.SUBCKT DLY4X1TS Y A VSS VDD
X0 net18 nmin VSS VSS LPNFET W=0.52U L=0.6U M=1 
X1 net21 net18 VSS VSS LPNFET W=0.52U L=0.6U M=1 
X2 net18 nmin VDD VDD LPPFET W=0.8U L=0.6U M=1 
X3 net21 net18 VDD VDD LPPFET W=0.8U L=0.6U M=1 
X4 VDD A nmin VDD LPPFET W=0.8U L=0.12U M=1 
X5 nmin A VSS VSS LPNFET W=0.52U L=0.12U M=1 
X6 VDD net21 Y VDD LPPFET W=0.64U L=0.12U M=1 
X7 Y net21 VSS VSS LPNFET W=0.24U L=0.12U M=1 
.ENDS DLY4X1TS 

**** 
*.SUBCKT DLY4X4TS Y A 
.SUBCKT DLY4X4TS Y A VSS VDD
X0 net18 nmin VSS VSS LPNFET W=0.58U L=0.56U M=1 
X1 net21 net18 VSS VSS LPNFET W=0.58U L=0.56U M=1 
X2 net18 nmin VDD VDD LPPFET W=0.8U L=0.56U M=1 
X3 net21 net18 VDD VDD LPPFET W=0.8U L=0.56U M=1 
X4 VDD A nmin VDD LPPFET W=0.8U L=0.12U M=1 
X5 nmin A VSS VSS LPNFET W=0.58U L=0.12U M=1 
X6 VDD net21 Y VDD LPPFET W=2.54U L=0.12U M=1 
X7 Y net21 VSS VSS LPNFET W=0.92U L=0.12U M=1 
.ENDS DLY4X4TS 

**** 
*.SUBCKT EDFFHQX1TS Q CK D E 
.SUBCKT EDFFHQX1TS Q CK D E VSS VDD
X0 VDD c hnet23 VDD LPPFET W=0.56U L=0.12U M=1 
X1 hnet23 nmin pm VDD LPPFET W=0.56U L=0.12U M=1 
X10 net98 c m VSS LPNFET W=0.46U L=0.12U M=1 
X11 hnet29 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X12 nmin nmen hnet29 VSS LPNFET W=0.2U L=0.12U M=1 
X13 hnet31 E nmin VDD LPPFET W=0.28U L=0.12U M=1 
X14 VDD s hnet31 VDD LPPFET W=0.28U L=0.12U M=1 
X15 hnet35 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X16 pm c hnet35 VSS LPNFET W=0.2U L=0.12U M=1 
X17 hnet37 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X18 VDD m hnet37 VDD LPPFET W=0.28U L=0.12U M=1 
X19 hnet41 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 hnet27 cn VSS VSS LPNFET W=0.4U L=0.12U M=1 
X20 net98 cn hnet41 VSS LPNFET W=0.2U L=0.12U M=1 
X21 hnet43 c net98 VDD LPPFET W=0.28U L=0.12U M=1 
X22 VDD s hnet43 VDD LPPFET W=0.28U L=0.12U M=1 
X23 VDD E nmen VDD LPPFET W=0.28U L=0.12U M=1 
X24 nmen E VSS VSS LPNFET W=0.2U L=0.12U M=1 
X25 VDD D net103 VDD LPPFET W=0.38U L=0.12U M=1 
X26 net103 D VSS VSS LPNFET W=0.28U L=0.12U M=1 
X27 VDD pm m VDD LPPFET W=0.92U L=0.12U M=1 
X28 m pm VSS VSS LPNFET W=0.48U L=0.12U M=1 
X29 VDD net98 s VDD LPPFET W=0.28U L=0.12U M=1 
X3 pm nmin hnet27 VSS LPNFET W=0.4U L=0.12U M=1 
X30 s net98 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X31 VDD net98 Q VDD LPPFET W=0.74U L=0.12U M=1 
X32 Q net98 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X33 VDD net113 c VDD LPPFET W=0.78U L=0.12U M=1 
X34 c net113 VSS VSS LPNFET W=0.28U L=0.12U M=1 
X35 VDD CK net113 VDD LPPFET W=0.28U L=0.12U M=1 
X36 net113 CK VSS VSS LPNFET W=0.28U L=0.12U M=1 
X4 net72 CK VDD VDD LPPFET W=0.7U L=0.12U M=1 
X5 cn c net72 VDD LPPFET W=0.52U L=0.12U M=1 
X6 nmin nmen net103 VDD LPPFET W=0.38U L=0.12U M=1 
X7 net98 cn m VDD LPPFET W=0.92U L=0.12U M=1 
X8 cn CK VSS VSS LPNFET W=0.2U L=0.12U M=1 
X9 nmin E net103 VSS LPNFET W=0.28U L=0.12U M=1 
.ENDS EDFFHQX1TS 

**** 
*.SUBCKT EDFFHQX2TS Q CK D E 
.SUBCKT EDFFHQX2TS Q CK D E VSS VDD
X0 VDD c hnet23 VDD LPPFET W=0.94U L=0.12U M=1 
X1 hnet23 nmin pm VDD LPPFET W=0.94U L=0.12U M=1 
X10 net98 c m VSS LPNFET W=0.74U L=0.12U M=1 
X11 hnet29 s VSS VSS LPNFET W=0.24U L=0.12U M=1 
X12 nmin nmen hnet29 VSS LPNFET W=0.24U L=0.12U M=1 
X13 hnet31 E nmin VDD LPPFET W=0.32U L=0.12U M=1 
X14 VDD s hnet31 VDD LPPFET W=0.32U L=0.12U M=1 
X15 hnet35 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X16 pm c hnet35 VSS LPNFET W=0.2U L=0.12U M=1 
X17 hnet37 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X18 VDD m hnet37 VDD LPPFET W=0.28U L=0.12U M=1 
X19 hnet41 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 hnet27 cn VSS VSS LPNFET W=0.68U L=0.12U M=1 
X20 net98 cn hnet41 VSS LPNFET W=0.2U L=0.12U M=1 
X21 hnet43 c net98 VDD LPPFET W=0.28U L=0.12U M=1 
X22 VDD s hnet43 VDD LPPFET W=0.28U L=0.12U M=1 
X23 VDD E nmen VDD LPPFET W=0.28U L=0.12U M=1 
X24 nmen E VSS VSS LPNFET W=0.2U L=0.12U M=1 
X25 VDD D net103 VDD LPPFET W=0.64U L=0.12U M=1 
X26 net103 D VSS VSS LPNFET W=0.46U L=0.12U M=1 
X27 VDD pm m VDD LPPFET W=1.3U L=0.12U M=1 
X28 m pm VSS VSS LPNFET W=0.8U L=0.12U M=1 
X29 VDD net98 s VDD LPPFET W=0.28U L=0.12U M=1 
X3 pm nmin hnet27 VSS LPNFET W=0.68U L=0.12U M=1 
X30 s net98 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X31 VDD net98 Q VDD LPPFET W=1.3U L=0.12U M=1 
X32 Q net98 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X33 VDD net113 c VDD LPPFET W=1.18U L=0.12U M=1 
X34 c net113 VSS VSS LPNFET W=0.42U L=0.12U M=1 
X35 VDD CK net113 VDD LPPFET W=0.32U L=0.12U M=1 
X36 net113 CK VSS VSS LPNFET W=0.32U L=0.12U M=1 
X4 net72 CK VDD VDD LPPFET W=0.9U L=0.12U M=1 
X5 cn c net72 VDD LPPFET W=0.68U L=0.12U M=1 
X6 nmin nmen net103 VDD LPPFET W=0.64U L=0.12U M=1 
X7 net98 cn m VDD LPPFET W=1.3U L=0.12U M=1 
X8 cn CK VSS VSS LPNFET W=0.26U L=0.12U M=1 
X9 nmin E net103 VSS LPNFET W=0.46U L=0.12U M=1 
.ENDS EDFFHQX2TS 

**** 
*.SUBCKT EDFFHQX4TS Q CK D E 
.SUBCKT EDFFHQX4TS Q CK D E VSS VDD
X0 hnet25 cn VSS VSS LPNFET W=0.66U L=0.12U M=1 
X1 pm nmin hnet25 VSS LPNFET W=0.66U L=0.12U M=1 
X10 net82 CK VDD VDD LPPFET W=0.76U L=0.12U M=1 
X11 cn c net82 VDD LPPFET W=0.64U L=0.12U M=1 
X12 nmin nmen net113 VDD LPPFET W=1.26U L=0.12U M=1 
X13 net108 cn m VDD LPPFET W=2.56U L=0.12U M=1 
X14 cn CK VSS VSS LPNFET W=0.48U L=0.12U M=1 
X15 nmin E net113 VSS LPNFET W=0.9U L=0.12U M=1 
X16 net108 c m VSS LPNFET W=1.38U L=0.12U M=1 
X17 hnet32 s VSS VSS LPNFET W=0.46U L=0.12U M=1 
X18 nmin nmen hnet32 VSS LPNFET W=0.46U L=0.12U M=1 
X19 hnet34 E nmin VDD LPPFET W=0.64U L=0.12U M=1 
X2 hnet21 cn VSS VSS LPNFET W=0.66U L=0.12U M=1 
X20 VDD s hnet34 VDD LPPFET W=0.64U L=0.12U M=1 
X21 hnet38 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X22 pm c hnet38 VSS LPNFET W=0.2U L=0.12U M=1 
X23 hnet40 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X24 VDD m hnet40 VDD LPPFET W=0.28U L=0.12U M=1 
X25 hnet44 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X26 net108 cn hnet44 VSS LPNFET W=0.2U L=0.12U M=1 
X27 hnet46 c net108 VDD LPPFET W=0.28U L=0.12U M=1 
X28 VDD s hnet46 VDD LPPFET W=0.28U L=0.12U M=1 
X29 VDD E nmen VDD LPPFET W=0.28U L=0.12U M=1 
X3 pm nmin hnet21 VSS LPNFET W=0.66U L=0.12U M=1 
X30 nmen E VSS VSS LPNFET W=0.2U L=0.12U M=1 
X31 VDD D net113 VDD LPPFET W=1.26U L=0.12U M=1 
X32 net113 D VSS VSS LPNFET W=0.9U L=0.12U M=1 
X33 VDD pm m VDD LPPFET W=2.76U L=0.12U M=1 
X34 m pm VSS VSS LPNFET W=1.58U L=0.12U M=1 
X35 VDD net108 s VDD LPPFET W=0.3U L=0.12U M=1 
X36 s net108 VSS VSS LPNFET W=0.22U L=0.12U M=1 
X37 VDD net108 Q VDD LPPFET W=2.6U L=0.12U M=1 
X38 Q net108 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X39 VDD net123 c VDD LPPFET W=2.02U L=0.12U M=1 
X4 VDD c hnet30 VDD LPPFET W=0.86U L=0.12U M=1 
X40 c net123 VSS VSS LPNFET W=0.72U L=0.12U M=1 
X41 VDD CK net123 VDD LPPFET W=0.54U L=0.12U M=1 
X42 net123 CK VSS VSS LPNFET W=0.54U L=0.12U M=1 
X5 hnet30 nmin pm VDD LPPFET W=0.86U L=0.12U M=1 
X6 VDD c hnet27 VDD LPPFET W=0.86U L=0.12U M=1 
X7 hnet27 nmin pm VDD LPPFET W=0.86U L=0.12U M=1 
X8 net76 CK VDD VDD LPPFET W=0.92U L=0.12U M=1 
X9 cn c net76 VDD LPPFET W=0.64U L=0.12U M=1 
.ENDS EDFFHQX4TS 

**** 
*.SUBCKT EDFFHQX8TS Q CK D E 
.SUBCKT EDFFHQX8TS Q CK D E VSS VDD
X0 hnet25 cn VSS VSS LPNFET W=0.66U L=0.12U M=1 
X1 pm nmin hnet25 VSS LPNFET W=0.66U L=0.12U M=1 
X10 net82 CK VDD VDD LPPFET W=0.76U L=0.12U M=1 
X11 cn c net82 VDD LPPFET W=0.64U L=0.12U M=1 
X12 nmin nmen net113 VDD LPPFET W=1.26U L=0.12U M=1 
X13 net108 cn m VDD LPPFET W=2.56U L=0.12U M=1 
X14 cn CK VSS VSS LPNFET W=0.48U L=0.12U M=1 
X15 nmin E net113 VSS LPNFET W=0.9U L=0.12U M=1 
X16 net108 c m VSS LPNFET W=1.38U L=0.12U M=1 
X17 hnet32 s VSS VSS LPNFET W=0.46U L=0.12U M=1 
X18 nmin nmen hnet32 VSS LPNFET W=0.46U L=0.12U M=1 
X19 hnet34 E nmin VDD LPPFET W=0.64U L=0.12U M=1 
X2 hnet21 cn VSS VSS LPNFET W=0.66U L=0.12U M=1 
X20 VDD s hnet34 VDD LPPFET W=0.64U L=0.12U M=1 
X21 hnet38 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X22 pm c hnet38 VSS LPNFET W=0.2U L=0.12U M=1 
X23 hnet40 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X24 VDD m hnet40 VDD LPPFET W=0.28U L=0.12U M=1 
X25 hnet44 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X26 net108 cn hnet44 VSS LPNFET W=0.2U L=0.12U M=1 
X27 hnet46 c net108 VDD LPPFET W=0.28U L=0.12U M=1 
X28 VDD s hnet46 VDD LPPFET W=0.28U L=0.12U M=1 
X29 VDD E nmen VDD LPPFET W=0.28U L=0.12U M=1 
X3 pm nmin hnet21 VSS LPNFET W=0.66U L=0.12U M=1 
X30 nmen E VSS VSS LPNFET W=0.2U L=0.12U M=1 
X31 VDD D net113 VDD LPPFET W=1.26U L=0.12U M=1 
X32 net113 D VSS VSS LPNFET W=0.9U L=0.12U M=1 
X33 VDD pm m VDD LPPFET W=2.76U L=0.12U M=1 
X34 m pm VSS VSS LPNFET W=1.58U L=0.12U M=1 
X35 VDD net108 s VDD LPPFET W=0.3U L=0.12U M=1 
X36 s net108 VSS VSS LPNFET W=0.22U L=0.12U M=1 
X37 VDD net108 Q VDD LPPFET W=5.2U L=0.12U M=1 
X38 Q net108 VSS VSS LPNFET W=3.68U L=0.12U M=1 
X39 VDD net123 c VDD LPPFET W=2.02U L=0.12U M=1 
X4 VDD c hnet30 VDD LPPFET W=0.86U L=0.12U M=1 
X40 c net123 VSS VSS LPNFET W=0.72U L=0.12U M=1 
X41 VDD CK net123 VDD LPPFET W=0.54U L=0.12U M=1 
X42 net123 CK VSS VSS LPNFET W=0.54U L=0.12U M=1 
X5 hnet30 nmin pm VDD LPPFET W=0.86U L=0.12U M=1 
X6 VDD c hnet27 VDD LPPFET W=0.86U L=0.12U M=1 
X7 hnet27 nmin pm VDD LPPFET W=0.86U L=0.12U M=1 
X8 net76 CK VDD VDD LPPFET W=0.92U L=0.12U M=1 
X9 cn c net76 VDD LPPFET W=0.64U L=0.12U M=1 
.ENDS EDFFHQX8TS 

**** 
*.SUBCKT EDFFTRX1TS Q QN CK D E RN 
.SUBCKT EDFFTRX1TS Q QN CK D E RN VSS VDD
X0 net72 RN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X1 net67 nmen net72 VSS LPNFET W=0.2U L=0.12U M=1 
X10 pm c net88 VDD LPPFET W=0.28U L=0.12U M=1 
X11 net88 RN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X12 VDD s net98 VDD LPPFET W=0.28U L=0.12U M=1 
X13 net98 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X14 VDD E nmen VDD LPPFET W=0.28U L=0.12U M=1 
X15 nmen E VSS VSS LPNFET W=0.2U L=0.12U M=1 
X16 VDD net98 Q VDD LPPFET W=0.64U L=0.12U M=1 
X17 Q net98 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X18 VDD s QN VDD LPPFET W=0.64U L=0.12U M=1 
X19 QN s VSS VSS LPNFET W=0.44U L=0.12U M=1 
X2 net76 s net67 VSS LPNFET W=0.2U L=0.12U M=1 
X20 VDD net115 s VDD LPPFET W=0.48U L=0.12U M=1 
X21 s net115 VSS VSS LPNFET W=0.34U L=0.12U M=1 
X22 VDD pm m VDD LPPFET W=0.28U L=0.12U M=1 
X23 m pm VSS VSS LPNFET W=0.2U L=0.12U M=1 
X24 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X25 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X26 VDD CK cn VDD LPPFET W=0.36U L=0.12U M=1 
X27 cn CK VSS VSS LPNFET W=0.26U L=0.12U M=1 
X28 hnet43 m VSS VSS LPNFET W=0.28U L=0.12U M=1 
X29 net115 c hnet43 VSS LPNFET W=0.28U L=0.12U M=1 
X3 net73 E net72 VSS LPNFET W=0.2U L=0.12U M=1 
X30 hnet45 cn net115 VDD LPPFET W=0.38U L=0.12U M=1 
X31 VDD m hnet45 VDD LPPFET W=0.38U L=0.12U M=1 
X32 hnet49 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X33 net115 cn hnet49 VSS LPNFET W=0.2U L=0.12U M=1 
X34 hnet51 c net115 VDD LPPFET W=0.28U L=0.12U M=1 
X35 VDD s hnet51 VDD LPPFET W=0.28U L=0.12U M=1 
X36 hnet55 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X37 pm c hnet55 VSS LPNFET W=0.2U L=0.12U M=1 
X38 hnet57 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X39 VDD m hnet57 VDD LPPFET W=0.28U L=0.12U M=1 
X4 net76 D net73 VSS LPNFET W=0.2U L=0.12U M=1 
X5 pm cn net76 VSS LPNFET W=0.2U L=0.12U M=1 
X6 net90 E VDD VDD LPPFET W=0.28U L=0.12U M=1 
X7 net87 nmen VDD VDD LPPFET W=0.28U L=0.12U M=1 
X8 net88 D net87 VDD LPPFET W=0.28U L=0.12U M=1 
X9 net88 s net90 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS EDFFTRX1TS 

**** 
*.SUBCKT EDFFTRX2TS Q QN CK D E RN 
.SUBCKT EDFFTRX2TS Q QN CK D E RN VSS VDD
X0 net72 RN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X1 net67 nmen net72 VSS LPNFET W=0.2U L=0.12U M=1 
X10 pm c net88 VDD LPPFET W=0.28U L=0.12U M=1 
X11 net88 RN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X12 VDD s net98 VDD LPPFET W=0.3U L=0.12U M=1 
X13 net98 s VSS VSS LPNFET W=0.22U L=0.12U M=1 
X14 VDD E nmen VDD LPPFET W=0.28U L=0.12U M=1 
X15 nmen E VSS VSS LPNFET W=0.2U L=0.12U M=1 
X16 VDD net98 Q VDD LPPFET W=1.28U L=0.12U M=1 
X17 Q net98 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X18 VDD s QN VDD LPPFET W=1.28U L=0.12U M=1 
X19 QN s VSS VSS LPNFET W=0.92U L=0.12U M=1 
X2 net76 s net67 VSS LPNFET W=0.2U L=0.12U M=1 
X20 VDD net115 s VDD LPPFET W=0.7U L=0.12U M=1 
X21 s net115 VSS VSS LPNFET W=0.5U L=0.12U M=1 
X22 VDD pm m VDD LPPFET W=0.28U L=0.12U M=1 
X23 m pm VSS VSS LPNFET W=0.2U L=0.12U M=1 
X24 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X25 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X26 VDD CK cn VDD LPPFET W=0.38U L=0.12U M=1 
X27 cn CK VSS VSS LPNFET W=0.28U L=0.12U M=1 
X28 hnet43 m VSS VSS LPNFET W=0.4U L=0.12U M=1 
X29 net115 c hnet43 VSS LPNFET W=0.4U L=0.12U M=1 
X3 net73 E net72 VSS LPNFET W=0.2U L=0.12U M=1 
X30 hnet45 cn net115 VDD LPPFET W=0.56U L=0.12U M=1 
X31 VDD m hnet45 VDD LPPFET W=0.56U L=0.12U M=1 
X32 hnet49 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X33 net115 cn hnet49 VSS LPNFET W=0.2U L=0.12U M=1 
X34 hnet51 c net115 VDD LPPFET W=0.28U L=0.12U M=1 
X35 VDD s hnet51 VDD LPPFET W=0.28U L=0.12U M=1 
X36 hnet55 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X37 pm c hnet55 VSS LPNFET W=0.2U L=0.12U M=1 
X38 hnet57 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X39 VDD m hnet57 VDD LPPFET W=0.28U L=0.12U M=1 
X4 net76 D net73 VSS LPNFET W=0.2U L=0.12U M=1 
X5 pm cn net76 VSS LPNFET W=0.2U L=0.12U M=1 
X6 net90 E VDD VDD LPPFET W=0.28U L=0.12U M=1 
X7 net87 nmen VDD VDD LPPFET W=0.28U L=0.12U M=1 
X8 net88 D net87 VDD LPPFET W=0.28U L=0.12U M=1 
X9 net88 s net90 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS EDFFTRX2TS 

**** 
*.SUBCKT EDFFTRX4TS Q QN CK D E RN 
.SUBCKT EDFFTRX4TS Q QN CK D E RN VSS VDD
X0 net73 RN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X1 net68 nmen net73 VSS LPNFET W=0.2U L=0.12U M=1 
X10 pm c net89 VDD LPPFET W=0.28U L=0.12U M=1 
X11 net89 RN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X12 VDD s net99 VDD LPPFET W=0.62U L=0.12U M=1 
X13 net99 s VSS VSS LPNFET W=0.44U L=0.12U M=1 
X14 VDD E nmen VDD LPPFET W=0.28U L=0.12U M=1 
X15 nmen E VSS VSS LPNFET W=0.2U L=0.12U M=1 
X16 VDD net99 Q VDD LPPFET W=2.56U L=0.12U M=1 
X17 Q net99 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X18 VDD s QN VDD LPPFET W=2.56U L=0.12U M=1 
X19 QN s VSS VSS LPNFET W=1.84U L=0.12U M=1 
X2 net77 s net68 VSS LPNFET W=0.2U L=0.12U M=1 
X20 VDD net116 s VDD LPPFET W=1.26U L=0.12U M=1 
X21 s net116 VSS VSS LPNFET W=0.9U L=0.12U M=1 
X22 VDD pm m VDD LPPFET W=0.36U L=0.12U M=1 
X23 m pm VSS VSS LPNFET W=0.26U L=0.12U M=1 
X24 VDD cn c VDD LPPFET W=0.34U L=0.12U M=1 
X25 c cn VSS VSS LPNFET W=0.24U L=0.12U M=1 
X26 VDD CK cn VDD LPPFET W=0.52U L=0.12U M=1 
X27 cn CK VSS VSS LPNFET W=0.38U L=0.12U M=1 
X28 hnet43 m VSS VSS LPNFET W=0.72U L=0.12U M=1 
X29 net116 c hnet43 VSS LPNFET W=0.72U L=0.12U M=1 
X3 net74 E net73 VSS LPNFET W=0.2U L=0.12U M=1 
X30 hnet45 cn net116 VDD LPPFET W=1U L=0.12U M=1 
X31 VDD m hnet45 VDD LPPFET W=1U L=0.12U M=1 
X32 hnet49 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X33 net116 cn hnet49 VSS LPNFET W=0.2U L=0.12U M=1 
X34 hnet51 c net116 VDD LPPFET W=0.28U L=0.12U M=1 
X35 VDD s hnet51 VDD LPPFET W=0.28U L=0.12U M=1 
X36 hnet55 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X37 pm c hnet55 VSS LPNFET W=0.2U L=0.12U M=1 
X38 hnet57 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X39 VDD m hnet57 VDD LPPFET W=0.28U L=0.12U M=1 
X4 net77 D net74 VSS LPNFET W=0.2U L=0.12U M=1 
X5 pm cn net77 VSS LPNFET W=0.2U L=0.12U M=1 
X6 net91 E VDD VDD LPPFET W=0.28U L=0.12U M=1 
X7 net88 nmen VDD VDD LPPFET W=0.28U L=0.12U M=1 
X8 net89 D net88 VDD LPPFET W=0.28U L=0.12U M=1 
X9 net89 s net91 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS EDFFTRX4TS 

**** 
*.SUBCKT EDFFTRXLTS Q QN CK D E RN 
.SUBCKT EDFFTRXLTS Q QN CK D E RN VSS VDD
X0 net73 RN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X1 net68 nmen net73 VSS LPNFET W=0.2U L=0.12U M=1 
X10 pm c net89 VDD LPPFET W=0.28U L=0.12U M=1 
X11 net89 RN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X12 VDD s net99 VDD LPPFET W=0.28U L=0.12U M=1 
X13 net99 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X14 VDD E nmen VDD LPPFET W=0.28U L=0.12U M=1 
X15 nmen E VSS VSS LPNFET W=0.2U L=0.12U M=1 
X16 VDD net99 Q VDD LPPFET W=0.34U L=0.12U M=1 
X17 Q net99 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X18 VDD s QN VDD LPPFET W=0.34U L=0.12U M=1 
X19 QN s VSS VSS LPNFET W=0.24U L=0.12U M=1 
X2 net77 s net68 VSS LPNFET W=0.2U L=0.12U M=1 
X20 VDD net116 s VDD LPPFET W=0.28U L=0.12U M=1 
X21 s net116 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X22 VDD pm m VDD LPPFET W=0.28U L=0.12U M=1 
X23 m pm VSS VSS LPNFET W=0.2U L=0.12U M=1 
X24 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X25 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X26 VDD CK cn VDD LPPFET W=0.34U L=0.12U M=1 
X27 cn CK VSS VSS LPNFET W=0.24U L=0.12U M=1 
X28 hnet43 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X29 net116 c hnet43 VSS LPNFET W=0.2U L=0.12U M=1 
X3 net74 E net73 VSS LPNFET W=0.2U L=0.12U M=1 
X30 hnet45 cn net116 VDD LPPFET W=0.28U L=0.12U M=1 
X31 VDD m hnet45 VDD LPPFET W=0.28U L=0.12U M=1 
X32 hnet49 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X33 net116 cn hnet49 VSS LPNFET W=0.2U L=0.12U M=1 
X34 hnet51 c net116 VDD LPPFET W=0.28U L=0.12U M=1 
X35 VDD s hnet51 VDD LPPFET W=0.28U L=0.12U M=1 
X36 hnet55 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X37 pm c hnet55 VSS LPNFET W=0.2U L=0.12U M=1 
X38 hnet57 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X39 VDD m hnet57 VDD LPPFET W=0.28U L=0.12U M=1 
X4 net77 D net74 VSS LPNFET W=0.2U L=0.12U M=1 
X5 pm cn net77 VSS LPNFET W=0.2U L=0.12U M=1 
X6 net91 E VDD VDD LPPFET W=0.28U L=0.12U M=1 
X7 net88 nmen VDD VDD LPPFET W=0.28U L=0.12U M=1 
X8 net89 D net88 VDD LPPFET W=0.28U L=0.12U M=1 
X9 net89 s net91 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS EDFFTRXLTS 

**** 
*.SUBCKT EDFFX1TS Q QN CK D E 
.SUBCKT EDFFX1TS Q QN CK D E VSS VDD
X0 net58 nmen VSS VSS LPNFET W=0.2U L=0.12U M=1 
X1 net67 s net58 VSS LPNFET W=0.2U L=0.12U M=1 
X10 VDD E nmen VDD LPPFET W=0.28U L=0.12U M=1 
X11 nmen E VSS VSS LPNFET W=0.2U L=0.12U M=1 
X12 VDD net101 Q VDD LPPFET W=0.64U L=0.12U M=1 
X13 Q net101 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X14 VDD s QN VDD LPPFET W=0.64U L=0.12U M=1 
X15 QN s VSS VSS LPNFET W=0.46U L=0.12U M=1 
X16 VDD net101 s VDD LPPFET W=0.28U L=0.12U M=1 
X17 s net101 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X18 VDD pm m VDD LPPFET W=0.28U L=0.12U M=1 
X19 m pm VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 net64 E VSS VSS LPNFET W=0.2U L=0.12U M=1 
X20 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X21 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X22 VDD CK cn VDD LPPFET W=0.3U L=0.12U M=1 
X23 cn CK VSS VSS LPNFET W=0.22U L=0.12U M=1 
X24 hnet38 m VSS VSS LPNFET W=0.22U L=0.12U M=1 
X25 net101 c hnet38 VSS LPNFET W=0.22U L=0.12U M=1 
X26 hnet40 cn net101 VDD LPPFET W=0.3U L=0.12U M=1 
X27 VDD m hnet40 VDD LPPFET W=0.3U L=0.12U M=1 
X28 hnet44 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X29 net101 cn hnet44 VSS LPNFET W=0.2U L=0.12U M=1 
X3 net67 D net64 VSS LPNFET W=0.2U L=0.12U M=1 
X30 hnet46 c net101 VDD LPPFET W=0.28U L=0.12U M=1 
X31 VDD s hnet46 VDD LPPFET W=0.28U L=0.12U M=1 
X32 hnet50 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X33 pm c hnet50 VSS LPNFET W=0.2U L=0.12U M=1 
X34 hnet52 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X35 VDD m hnet52 VDD LPPFET W=0.28U L=0.12U M=1 
X4 pm cn net67 VSS LPNFET W=0.2U L=0.12U M=1 
X5 net81 E VDD VDD LPPFET W=0.28U L=0.12U M=1 
X6 net78 nmen VDD VDD LPPFET W=0.28U L=0.12U M=1 
X7 net79 D net78 VDD LPPFET W=0.28U L=0.12U M=1 
X8 net79 s net81 VDD LPPFET W=0.28U L=0.12U M=1 
X9 pm c net79 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS EDFFX1TS 

**** 
*.SUBCKT EDFFX2TS Q QN CK D E 
.SUBCKT EDFFX2TS Q QN CK D E VSS VDD
X0 net58 nmen VSS VSS LPNFET W=0.2U L=0.12U M=1 
X1 net67 s net58 VSS LPNFET W=0.2U L=0.12U M=1 
X10 VDD E nmen VDD LPPFET W=0.28U L=0.12U M=1 
X11 nmen E VSS VSS LPNFET W=0.2U L=0.12U M=1 
X12 VDD net101 Q VDD LPPFET W=1.28U L=0.12U M=1 
X13 Q net101 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X14 VDD s QN VDD LPPFET W=1.2U L=0.12U M=1 
X15 QN s VSS VSS LPNFET W=0.92U L=0.12U M=1 
X16 VDD net101 s VDD LPPFET W=0.28U L=0.12U M=1 
X17 s net101 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X18 VDD pm m VDD LPPFET W=0.28U L=0.12U M=1 
X19 m pm VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 net64 E VSS VSS LPNFET W=0.2U L=0.12U M=1 
X20 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X21 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X22 VDD CK cn VDD LPPFET W=0.36U L=0.12U M=1 
X23 cn CK VSS VSS LPNFET W=0.26U L=0.12U M=1 
X24 hnet38 m VSS VSS LPNFET W=0.4U L=0.12U M=1 
X25 net101 c hnet38 VSS LPNFET W=0.4U L=0.12U M=1 
X26 hnet40 cn net101 VDD LPPFET W=0.52U L=0.12U M=1 
X27 VDD m hnet40 VDD LPPFET W=0.52U L=0.12U M=1 
X28 hnet44 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X29 net101 cn hnet44 VSS LPNFET W=0.2U L=0.12U M=1 
X3 net67 D net64 VSS LPNFET W=0.2U L=0.12U M=1 
X30 hnet46 c net101 VDD LPPFET W=0.28U L=0.12U M=1 
X31 VDD s hnet46 VDD LPPFET W=0.28U L=0.12U M=1 
X32 hnet50 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X33 pm c hnet50 VSS LPNFET W=0.2U L=0.12U M=1 
X34 hnet52 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X35 VDD m hnet52 VDD LPPFET W=0.28U L=0.12U M=1 
X4 pm cn net67 VSS LPNFET W=0.2U L=0.12U M=1 
X5 net81 E VDD VDD LPPFET W=0.28U L=0.12U M=1 
X6 net78 nmen VDD VDD LPPFET W=0.28U L=0.12U M=1 
X7 net79 D net78 VDD LPPFET W=0.28U L=0.12U M=1 
X8 net79 s net81 VDD LPPFET W=0.28U L=0.12U M=1 
X9 pm c net79 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS EDFFX2TS 

**** 
*.SUBCKT EDFFX4TS Q QN CK D E 
.SUBCKT EDFFX4TS Q QN CK D E VSS VDD
X0 hnet24 m VSS VSS LPNFET W=0.38U L=0.12U M=1 
X1 hnet25 m VSS VSS LPNFET W=0.38U L=0.12U M=1 
X10 net67 E VSS VSS LPNFET W=0.2U L=0.12U M=1 
X11 net70 D net67 VSS LPNFET W=0.2U L=0.12U M=1 
X12 pm cn net70 VSS LPNFET W=0.2U L=0.12U M=1 
X13 net84 E VDD VDD LPPFET W=0.28U L=0.12U M=1 
X14 net81 nmen VDD VDD LPPFET W=0.28U L=0.12U M=1 
X15 net82 D net81 VDD LPPFET W=0.28U L=0.12U M=1 
X16 net82 s net84 VDD LPPFET W=0.28U L=0.12U M=1 
X17 pm c net82 VDD LPPFET W=0.28U L=0.12U M=1 
X18 VDD E nmen VDD LPPFET W=0.28U L=0.12U M=1 
X19 nmen E VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 net56 c hnet24 VSS LPNFET W=0.38U L=0.12U M=1 
X20 VDD net56 Q VDD LPPFET W=2.56U L=0.12U M=1 
X21 Q net56 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X22 VDD s QN VDD LPPFET W=2.56U L=0.12U M=1 
X23 QN s VSS VSS LPNFET W=1.84U L=0.12U M=1 
X24 VDD net56 s VDD LPPFET W=0.52U L=0.12U M=1 
X25 s net56 VSS VSS LPNFET W=0.38U L=0.12U M=1 
X26 VDD pm m VDD LPPFET W=0.28U L=0.12U M=1 
X27 m pm VSS VSS LPNFET W=0.2U L=0.12U M=1 
X28 VDD cn c VDD LPPFET W=0.34U L=0.12U M=1 
X29 c cn VSS VSS LPNFET W=0.24U L=0.12U M=1 
X3 net56 c hnet25 VSS LPNFET W=0.38U L=0.12U M=1 
X30 VDD CK cn VDD LPPFET W=0.5U L=0.12U M=1 
X31 cn CK VSS VSS LPNFET W=0.36U L=0.12U M=1 
X32 hnet46 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X33 net56 cn hnet46 VSS LPNFET W=0.2U L=0.12U M=1 
X34 hnet48 c net56 VDD LPPFET W=0.28U L=0.12U M=1 
X35 VDD s hnet48 VDD LPPFET W=0.28U L=0.12U M=1 
X36 hnet52 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X37 pm c hnet52 VSS LPNFET W=0.2U L=0.12U M=1 
X38 hnet54 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X39 VDD m hnet54 VDD LPPFET W=0.28U L=0.12U M=1 
X4 hnet30 cn net56 VDD LPPFET W=0.54U L=0.12U M=1 
X5 hnet28 cn net56 VDD LPPFET W=0.54U L=0.12U M=1 
X6 VDD m hnet30 VDD LPPFET W=0.54U L=0.12U M=1 
X7 VDD m hnet28 VDD LPPFET W=0.54U L=0.12U M=1 
X8 net61 nmen VSS VSS LPNFET W=0.2U L=0.12U M=1 
X9 net70 s net61 VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS EDFFX4TS 

**** 
*.SUBCKT EDFFXLTS Q QN CK D E 
.SUBCKT EDFFXLTS Q QN CK D E VSS VDD
X0 net58 nmen VSS VSS LPNFET W=0.2U L=0.12U M=1 
X1 net67 s net58 VSS LPNFET W=0.2U L=0.12U M=1 
X10 VDD E nmen VDD LPPFET W=0.28U L=0.12U M=1 
X11 nmen E VSS VSS LPNFET W=0.2U L=0.12U M=1 
X12 VDD net101 Q VDD LPPFET W=0.34U L=0.12U M=1 
X13 Q net101 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X14 VDD s QN VDD LPPFET W=0.34U L=0.12U M=1 
X15 QN s VSS VSS LPNFET W=0.24U L=0.12U M=1 
X16 VDD net101 s VDD LPPFET W=0.28U L=0.12U M=1 
X17 s net101 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X18 VDD pm m VDD LPPFET W=0.28U L=0.12U M=1 
X19 m pm VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 net64 E VSS VSS LPNFET W=0.2U L=0.12U M=1 
X20 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X21 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X22 VDD CK cn VDD LPPFET W=0.3U L=0.12U M=1 
X23 cn CK VSS VSS LPNFET W=0.22U L=0.12U M=1 
X24 hnet38 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X25 net101 c hnet38 VSS LPNFET W=0.2U L=0.12U M=1 
X26 hnet40 cn net101 VDD LPPFET W=0.28U L=0.12U M=1 
X27 VDD m hnet40 VDD LPPFET W=0.28U L=0.12U M=1 
X28 hnet44 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X29 net101 cn hnet44 VSS LPNFET W=0.2U L=0.12U M=1 
X3 net67 D net64 VSS LPNFET W=0.2U L=0.12U M=1 
X30 hnet46 c net101 VDD LPPFET W=0.28U L=0.12U M=1 
X31 VDD s hnet46 VDD LPPFET W=0.28U L=0.12U M=1 
X32 hnet50 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X33 pm c hnet50 VSS LPNFET W=0.2U L=0.12U M=1 
X34 hnet52 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X35 VDD m hnet52 VDD LPPFET W=0.28U L=0.12U M=1 
X4 pm cn net67 VSS LPNFET W=0.2U L=0.12U M=1 
X5 net81 E VDD VDD LPPFET W=0.28U L=0.12U M=1 
X6 net78 nmen VDD VDD LPPFET W=0.28U L=0.12U M=1 
X7 net79 D net78 VDD LPPFET W=0.28U L=0.12U M=1 
X8 net79 s net81 VDD LPPFET W=0.28U L=0.12U M=1 
X9 pm c net79 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS EDFFXLTS 

**** 
*.SUBCKT HOLDX1TS Y 
.SUBCKT HOLDX1TS Y VSS VDD
X0 Y nmio net11 VSS LPNFET W=0.2U L=0.12U M=1 
X1 net11 nmio VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 Y nmio VDD VDD LPPFET W=0.28U L=0.12U M=1 
X3 VDD Y nmio VDD LPPFET W=0.28U L=0.12U M=1 
X4 nmio Y VSS VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS HOLDX1TS 

**** 
*.SUBCKT INVX12TS Y A 
.SUBCKT INVX12TS Y A VSS VDD
X0 VDD A Y VDD LPPFET W=7.54U L=0.12U M=1 
X1 Y A VSS VSS LPNFET W=5.26U L=0.12U M=1 
.ENDS INVX12TS 

**** 
*.SUBCKT INVX16TS Y A 
.SUBCKT INVX16TS Y A VSS VDD
X0 VDD A Y VDD LPPFET W=10.2U L=0.12U M=1 
X1 Y A VSS VSS LPNFET W=7.1U L=0.12U M=1 
.ENDS INVX16TS 

**** 
*.SUBCKT INVX1TS Y A 
.SUBCKT INVX1TS Y A VSS VDD
X0 VDD A Y VDD LPPFET W=0.64U L=0.12U M=1 
X1 Y A VSS VSS LPNFET W=0.46U L=0.12U M=1 
.ENDS INVX1TS 

**** 
*.SUBCKT INVX20TS Y A 
.SUBCKT INVX20TS Y A VSS VDD
X0 VDD A Y VDD LPPFET W=12.5U L=0.12U M=1 
X1 Y A VSS VSS LPNFET W=8.68U L=0.12U M=1 
.ENDS INVX20TS 

**** 
*.SUBCKT INVX2TS Y A 
.SUBCKT INVX2TS Y A VSS VDD
X0 VDD A Y VDD LPPFET W=1.28U L=0.12U M=1 
X1 Y A VSS VSS LPNFET W=0.92U L=0.12U M=1 
.ENDS INVX2TS 

**** 
*.SUBCKT INVX3TS Y A 
.SUBCKT INVX3TS Y A VSS VDD
X0 VDD A Y VDD LPPFET W=1.9U L=0.12U M=1 
X1 Y A VSS VSS LPNFET W=1.32U L=0.12U M=1 
.ENDS INVX3TS 

**** 
*.SUBCKT INVX4TS Y A 
.SUBCKT INVX4TS Y A VSS VDD
X0 VDD A Y VDD LPPFET W=2.34U L=0.12U M=1 
X1 Y A VSS VSS LPNFET W=1.7U L=0.12U M=1 
.ENDS INVX4TS 

**** 
*.SUBCKT INVX6TS Y A 
.SUBCKT INVX6TS Y A VSS VDD
X0 VDD A Y VDD LPPFET W=3.76U L=0.12U M=1 
X1 Y A VSS VSS LPNFET W=2.56U L=0.12U M=1 
.ENDS INVX6TS 

**** 
*.SUBCKT INVX8TS Y A 
.SUBCKT INVX8TS Y A VSS VDD
X0 VDD A Y VDD LPPFET W=4.96U L=0.12U M=1 
X1 Y A VSS VSS LPNFET W=3.42U L=0.12U M=1 
.ENDS INVX8TS 

**** 
*.SUBCKT INVXLTS Y A 
.SUBCKT INVXLTS Y A VSS VDD
X0 VDD A Y VDD LPPFET W=0.34U L=0.12U M=1 
X1 Y A VSS VSS LPNFET W=0.24U L=0.12U M=1 
.ENDS INVXLTS 

**** 
*.SUBCKT MDFFHQX1TS Q CK D0 D1 S0 
.SUBCKT MDFFHQX1TS Q CK D0 D1 S0 VSS VDD
X0 VDD c hnet25 VDD LPPFET W=0.58U L=0.12U M=1 
X1 hnet25 net87 pm VDD LPPFET W=0.58U L=0.12U M=1 
X10 net87 nmsel nmin0 VSS LPNFET W=0.28U L=0.12U M=1 
X11 net87 S0 nmin1 VSS LPNFET W=0.3U L=0.12U M=1 
X12 net99 c m VSS LPNFET W=0.48U L=0.12U M=1 
X13 hnet31 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X14 pm c hnet31 VSS LPNFET W=0.2U L=0.12U M=1 
X15 hnet33 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X16 VDD m hnet33 VDD LPPFET W=0.28U L=0.12U M=1 
X17 hnet37 s VSS VSS LPNFET W=0.18U L=0.12U M=1 
X18 net99 cn hnet37 VSS LPNFET W=0.18U L=0.12U M=1 
X19 hnet39 c net99 VDD LPPFET W=0.28U L=0.12U M=1 
X2 hnet29 cn VSS VSS LPNFET W=0.42U L=0.12U M=1 
X20 VDD s hnet39 VDD LPPFET W=0.28U L=0.12U M=1 
X21 VDD D0 nmin0 VDD LPPFET W=0.38U L=0.12U M=1 
X22 nmin0 D0 VSS VSS LPNFET W=0.28U L=0.12U M=1 
X23 VDD D1 nmin1 VDD LPPFET W=0.38U L=0.12U M=1 
X24 nmin1 D1 VSS VSS LPNFET W=0.3U L=0.12U M=1 
X25 VDD S0 nmsel VDD LPPFET W=0.48U L=0.12U M=1 
X26 nmsel S0 VSS VSS LPNFET W=0.34U L=0.12U M=1 
X27 VDD pm m VDD LPPFET W=0.96U L=0.12U M=1 
X28 m pm VSS VSS LPNFET W=0.5U L=0.12U M=1 
X29 VDD net99 s VDD LPPFET W=0.28U L=0.12U M=1 
X3 pm net87 hnet29 VSS LPNFET W=0.42U L=0.12U M=1 
X30 s net99 VSS VSS LPNFET W=0.18U L=0.12U M=1 
X31 VDD net99 Q VDD LPPFET W=0.74U L=0.12U M=1 
X32 Q net99 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X33 VDD net116 c VDD LPPFET W=0.84U L=0.12U M=1 
X34 c net116 VSS VSS LPNFET W=0.3U L=0.12U M=1 
X35 VDD CK net116 VDD LPPFET W=0.28U L=0.12U M=1 
X36 net116 CK VSS VSS LPNFET W=0.28U L=0.12U M=1 
X4 net71 CK VDD VDD LPPFET W=0.7U L=0.12U M=1 
X5 cn c net71 VDD LPPFET W=0.52U L=0.12U M=1 
X6 net87 S0 nmin0 VDD LPPFET W=0.38U L=0.12U M=1 
X7 net87 nmsel nmin1 VDD LPPFET W=0.38U L=0.12U M=1 
X8 net99 cn m VDD LPPFET W=0.96U L=0.12U M=1 
X9 cn CK VSS VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS MDFFHQX1TS 

**** 
*.SUBCKT MDFFHQX2TS Q CK D0 D1 S0 
.SUBCKT MDFFHQX2TS Q CK D0 D1 S0 VSS VDD
X0 VDD c hnet25 VDD LPPFET W=1U L=0.12U M=1 
X1 hnet25 net87 pm VDD LPPFET W=1U L=0.12U M=1 
X10 net87 nmsel nmin0 VSS LPNFET W=0.48U L=0.12U M=1 
X11 net87 S0 nmin1 VSS LPNFET W=0.5U L=0.12U M=1 
X12 net99 c m VSS LPNFET W=0.72U L=0.12U M=1 
X13 hnet31 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X14 pm c hnet31 VSS LPNFET W=0.2U L=0.12U M=1 
X15 hnet33 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X16 VDD m hnet33 VDD LPPFET W=0.28U L=0.12U M=1 
X17 hnet37 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X18 net99 cn hnet37 VSS LPNFET W=0.2U L=0.12U M=1 
X19 hnet39 c net99 VDD LPPFET W=0.28U L=0.12U M=1 
X2 hnet29 cn VSS VSS LPNFET W=0.66U L=0.12U M=1 
X20 VDD s hnet39 VDD LPPFET W=0.28U L=0.12U M=1 
X21 VDD D0 nmin0 VDD LPPFET W=0.68U L=0.12U M=1 
X22 nmin0 D0 VSS VSS LPNFET W=0.48U L=0.12U M=1 
X23 VDD D1 nmin1 VDD LPPFET W=0.68U L=0.12U M=1 
X24 nmin1 D1 VSS VSS LPNFET W=0.5U L=0.12U M=1 
X25 VDD S0 nmsel VDD LPPFET W=0.84U L=0.12U M=1 
X26 nmsel S0 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X27 VDD pm m VDD LPPFET W=1.48U L=0.12U M=1 
X28 m pm VSS VSS LPNFET W=0.72U L=0.12U M=1 
X29 VDD net99 s VDD LPPFET W=0.28U L=0.12U M=1 
X3 pm net87 hnet29 VSS LPNFET W=0.66U L=0.12U M=1 
X30 s net99 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X31 VDD net99 Q VDD LPPFET W=1.56U L=0.12U M=1 
X32 Q net99 VSS VSS LPNFET W=0.76U L=0.12U M=1 
X33 VDD net116 c VDD LPPFET W=1.2U L=0.12U M=1 
X34 c net116 VSS VSS LPNFET W=0.42U L=0.12U M=1 
X35 VDD CK net116 VDD LPPFET W=0.32U L=0.12U M=1 
X36 net116 CK VSS VSS LPNFET W=0.28U L=0.12U M=1 
X4 net71 CK VDD VDD LPPFET W=0.84U L=0.12U M=1 
X5 cn c net71 VDD LPPFET W=0.68U L=0.12U M=1 
X6 net87 S0 nmin0 VDD LPPFET W=0.68U L=0.12U M=1 
X7 net87 nmsel nmin1 VDD LPPFET W=0.68U L=0.12U M=1 
X8 net99 cn m VDD LPPFET W=1.36U L=0.12U M=1 
X9 cn CK VSS VSS LPNFET W=0.26U L=0.12U M=1 
.ENDS MDFFHQX2TS 

**** 
*.SUBCKT MDFFHQX4TS Q CK D0 D1 S0 
.SUBCKT MDFFHQX4TS Q CK D0 D1 S0 VSS VDD
X0 hnet27 cn VSS VSS LPNFET W=0.66U L=0.12U M=1 
X1 pm net93 hnet27 VSS LPNFET W=0.66U L=0.12U M=1 
X10 net77 CK VDD VDD LPPFET W=0.84U L=0.12U M=1 
X11 cn c net77 VDD LPPFET W=0.64U L=0.12U M=1 
X12 net93 S0 nmin0 VDD LPPFET W=1.22U L=0.12U M=1 
X13 net93 nmsel nmin1 VDD LPPFET W=1.22U L=0.12U M=1 
X14 net105 cn m VDD LPPFET W=2.72U L=0.12U M=1 
X15 cn CK VSS VSS LPNFET W=0.48U L=0.12U M=1 
X16 net93 nmsel nmin0 VSS LPNFET W=0.88U L=0.12U M=1 
X17 net93 S0 nmin1 VSS LPNFET W=0.88U L=0.12U M=1 
X18 net105 c m VSS LPNFET W=1.5U L=0.12U M=1 
X19 hnet34 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 hnet23 cn VSS VSS LPNFET W=0.66U L=0.12U M=1 
X20 pm c hnet34 VSS LPNFET W=0.2U L=0.12U M=1 
X21 hnet36 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X22 VDD m hnet36 VDD LPPFET W=0.28U L=0.12U M=1 
X23 hnet40 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X24 net105 cn hnet40 VSS LPNFET W=0.2U L=0.12U M=1 
X25 hnet42 c net105 VDD LPPFET W=0.28U L=0.12U M=1 
X26 VDD s hnet42 VDD LPPFET W=0.28U L=0.12U M=1 
X27 VDD D0 nmin0 VDD LPPFET W=1.22U L=0.12U M=1 
X28 nmin0 D0 VSS VSS LPNFET W=0.88U L=0.12U M=1 
X29 VDD D1 nmin1 VDD LPPFET W=1.22U L=0.12U M=1 
X3 pm net93 hnet23 VSS LPNFET W=0.66U L=0.12U M=1 
X30 nmin1 D1 VSS VSS LPNFET W=0.88U L=0.12U M=1 
X31 VDD S0 nmsel VDD LPPFET W=1.5U L=0.12U M=1 
X32 nmsel S0 VSS VSS LPNFET W=1.08U L=0.12U M=1 
X33 VDD pm m VDD LPPFET W=2.72U L=0.12U M=1 
X34 m pm VSS VSS LPNFET W=1.32U L=0.12U M=1 
X35 VDD net105 s VDD LPPFET W=0.28U L=0.12U M=1 
X36 s net105 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X37 VDD net105 Q VDD LPPFET W=2.6U L=0.12U M=1 
X38 Q net105 VSS VSS LPNFET W=1.82U L=0.12U M=1 
X39 VDD net122 c VDD LPPFET W=2.02U L=0.12U M=1 
X4 VDD c hnet32 VDD LPPFET W=0.9U L=0.12U M=1 
X40 c net122 VSS VSS LPNFET W=0.72U L=0.12U M=1 
X41 VDD CK net122 VDD LPPFET W=0.54U L=0.12U M=1 
X42 net122 CK VSS VSS LPNFET W=0.54U L=0.12U M=1 
X5 hnet32 net93 pm VDD LPPFET W=0.9U L=0.12U M=1 
X6 VDD c hnet29 VDD LPPFET W=0.9U L=0.12U M=1 
X7 hnet29 net93 pm VDD LPPFET W=0.9U L=0.12U M=1 
X8 net71 CK VDD VDD LPPFET W=0.84U L=0.12U M=1 
X9 cn c net71 VDD LPPFET W=0.64U L=0.12U M=1 
.ENDS MDFFHQX4TS 

**** 
*.SUBCKT MDFFHQX8TS Q CK D0 D1 S0 
.SUBCKT MDFFHQX8TS Q CK D0 D1 S0 VSS VDD
X0 hnet27 cn VSS VSS LPNFET W=0.66U L=0.12U M=1 
X1 pm net93 hnet27 VSS LPNFET W=0.66U L=0.12U M=1 
X10 net77 CK VDD VDD LPPFET W=0.84U L=0.12U M=1 
X11 cn c net77 VDD LPPFET W=0.64U L=0.12U M=1 
X12 net93 S0 nmin0 VDD LPPFET W=1.22U L=0.12U M=1 
X13 net93 nmsel nmin1 VDD LPPFET W=1.22U L=0.12U M=1 
X14 net105 cn m VDD LPPFET W=2.72U L=0.12U M=1 
X15 cn CK VSS VSS LPNFET W=0.48U L=0.12U M=1 
X16 net93 nmsel nmin0 VSS LPNFET W=0.88U L=0.12U M=1 
X17 net93 S0 nmin1 VSS LPNFET W=0.88U L=0.12U M=1 
X18 net105 c m VSS LPNFET W=1.5U L=0.12U M=1 
X19 hnet34 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 hnet23 cn VSS VSS LPNFET W=0.66U L=0.12U M=1 
X20 pm c hnet34 VSS LPNFET W=0.2U L=0.12U M=1 
X21 hnet36 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X22 VDD m hnet36 VDD LPPFET W=0.28U L=0.12U M=1 
X23 hnet40 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X24 net105 cn hnet40 VSS LPNFET W=0.2U L=0.12U M=1 
X25 hnet42 c net105 VDD LPPFET W=0.28U L=0.12U M=1 
X26 VDD s hnet42 VDD LPPFET W=0.28U L=0.12U M=1 
X27 VDD D0 nmin0 VDD LPPFET W=1.22U L=0.12U M=1 
X28 nmin0 D0 VSS VSS LPNFET W=0.88U L=0.12U M=1 
X29 VDD D1 nmin1 VDD LPPFET W=1.22U L=0.12U M=1 
X3 pm net93 hnet23 VSS LPNFET W=0.66U L=0.12U M=1 
X30 nmin1 D1 VSS VSS LPNFET W=0.88U L=0.12U M=1 
X31 VDD S0 nmsel VDD LPPFET W=1.5U L=0.12U M=1 
X32 nmsel S0 VSS VSS LPNFET W=1.08U L=0.12U M=1 
X33 VDD pm m VDD LPPFET W=2.72U L=0.12U M=1 
X34 m pm VSS VSS LPNFET W=1.32U L=0.12U M=1 
X35 VDD net105 s VDD LPPFET W=0.28U L=0.12U M=1 
X36 s net105 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X37 VDD net105 Q VDD LPPFET W=5.2U L=0.12U M=1 
X38 Q net105 VSS VSS LPNFET W=3.64U L=0.12U M=1 
X39 VDD net122 c VDD LPPFET W=2.02U L=0.12U M=1 
X4 VDD c hnet32 VDD LPPFET W=0.9U L=0.12U M=1 
X40 c net122 VSS VSS LPNFET W=0.72U L=0.12U M=1 
X41 VDD CK net122 VDD LPPFET W=0.54U L=0.12U M=1 
X42 net122 CK VSS VSS LPNFET W=0.54U L=0.12U M=1 
X5 hnet32 net93 pm VDD LPPFET W=0.9U L=0.12U M=1 
X6 VDD c hnet29 VDD LPPFET W=0.9U L=0.12U M=1 
X7 hnet29 net93 pm VDD LPPFET W=0.9U L=0.12U M=1 
X8 net71 CK VDD VDD LPPFET W=0.84U L=0.12U M=1 
X9 cn c net71 VDD LPPFET W=0.64U L=0.12U M=1 
.ENDS MDFFHQX8TS 

**** 
*.SUBCKT MX2X1TS Y A B S0 
.SUBCKT MX2X1TS Y A B S0 VSS VDD
X0 net25 nmsel nmin0 VSS LPNFET W=0.36U L=0.12U M=1 
X1 net25 S0 nmin1 VSS LPNFET W=0.36U L=0.12U M=1 
X10 VDD S0 nmsel VDD LPPFET W=0.28U L=0.12U M=1 
X11 nmsel S0 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 net25 S0 nmin0 VDD LPPFET W=0.5U L=0.12U M=1 
X3 net25 nmsel nmin1 VDD LPPFET W=0.5U L=0.12U M=1 
X4 VDD net25 Y VDD LPPFET W=0.64U L=0.12U M=1 
X5 Y net25 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X6 VDD A nmin0 VDD LPPFET W=0.5U L=0.12U M=1 
X7 nmin0 A VSS VSS LPNFET W=0.36U L=0.12U M=1 
X8 VDD B nmin1 VDD LPPFET W=0.5U L=0.12U M=1 
X9 nmin1 B VSS VSS LPNFET W=0.36U L=0.12U M=1 
.ENDS MX2X1TS 

**** 
*.SUBCKT MX2X2TS Y A B S0 
.SUBCKT MX2X2TS Y A B S0 VSS VDD
X0 net25 nmsel nmin0 VSS LPNFET W=0.74U L=0.12U M=1 
X1 net25 S0 nmin1 VSS LPNFET W=0.74U L=0.12U M=1 
X10 VDD S0 nmsel VDD LPPFET W=0.42U L=0.12U M=1 
X11 nmsel S0 VSS VSS LPNFET W=0.3U L=0.12U M=1 
X2 net25 S0 nmin0 VDD LPPFET W=0.98U L=0.12U M=1 
X3 net25 nmsel nmin1 VDD LPPFET W=0.98U L=0.12U M=1 
X4 VDD net25 Y VDD LPPFET W=1.28U L=0.12U M=1 
X5 Y net25 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X6 VDD A nmin0 VDD LPPFET W=0.98U L=0.12U M=1 
X7 nmin0 A VSS VSS LPNFET W=0.74U L=0.12U M=1 
X8 VDD B nmin1 VDD LPPFET W=0.98U L=0.12U M=1 
X9 nmin1 B VSS VSS LPNFET W=0.74U L=0.12U M=1 
.ENDS MX2X2TS 

**** 
*.SUBCKT MX2X4TS Y A B S0 
.SUBCKT MX2X4TS Y A B S0 VSS VDD
X0 net25 nmsel nmin0 VSS LPNFET W=0.82U L=0.12U M=1 
X1 net25 S0 nmin1 VSS LPNFET W=0.82U L=0.12U M=1 
X10 VDD S0 nmsel VDD LPPFET W=0.5U L=0.12U M=1 
X11 nmsel S0 VSS VSS LPNFET W=0.36U L=0.12U M=1 
X2 net25 S0 nmin0 VDD LPPFET W=1.28U L=0.12U M=1 
X3 net25 nmsel nmin1 VDD LPPFET W=1.28U L=0.12U M=1 
X4 VDD net25 Y VDD LPPFET W=2.56U L=0.12U M=1 
X5 Y net25 VSS VSS LPNFET W=1.64U L=0.12U M=1 
X6 VDD A nmin0 VDD LPPFET W=1.28U L=0.12U M=1 
X7 nmin0 A VSS VSS LPNFET W=0.82U L=0.12U M=1 
X8 VDD B nmin1 VDD LPPFET W=1.28U L=0.12U M=1 
X9 nmin1 B VSS VSS LPNFET W=0.82U L=0.12U M=1 
.ENDS MX2X4TS 

**** 
*.SUBCKT MX2X6TS Y A B S0 
.SUBCKT MX2X6TS Y A B S0 VSS VDD
X0 net25 nmsel nmin0 VSS LPNFET W=0.8U L=0.12U M=1 
X1 net25 S0 nmin1 VSS LPNFET W=0.8U L=0.12U M=1 
X10 VDD S0 nmsel VDD LPPFET W=0.5U L=0.12U M=1 
X11 nmsel S0 VSS VSS LPNFET W=0.36U L=0.12U M=1 
X2 net25 S0 nmin0 VDD LPPFET W=1.28U L=0.12U M=1 
X3 net25 nmsel nmin1 VDD LPPFET W=1.28U L=0.12U M=1 
X4 VDD net25 Y VDD LPPFET W=3.84U L=0.12U M=1 
X5 Y net25 VSS VSS LPNFET W=2.76U L=0.12U M=1 
X6 VDD A nmin0 VDD LPPFET W=1.28U L=0.12U M=1 
X7 nmin0 A VSS VSS LPNFET W=0.92U L=0.12U M=1 
X8 VDD B nmin1 VDD LPPFET W=1.28U L=0.12U M=1 
X9 nmin1 B VSS VSS LPNFET W=0.92U L=0.12U M=1 
.ENDS MX2X6TS 

**** 
*.SUBCKT MX2X8TS Y A B S0 
.SUBCKT MX2X8TS Y A B S0 VSS VDD
X0 net25 nmsel nmin0 VSS LPNFET W=0.76U L=0.12U M=1 
X1 net25 S0 nmin1 VSS LPNFET W=0.76U L=0.12U M=1 
X10 VDD S0 nmsel VDD LPPFET W=0.5U L=0.12U M=1 
X11 nmsel S0 VSS VSS LPNFET W=0.36U L=0.12U M=1 
X2 net25 S0 nmin0 VDD LPPFET W=1.24U L=0.12U M=1 
X3 net25 nmsel nmin1 VDD LPPFET W=1.24U L=0.12U M=1 
X4 VDD net25 Y VDD LPPFET W=5.12U L=0.12U M=1 
X5 Y net25 VSS VSS LPNFET W=3.32U L=0.12U M=1 
X6 VDD A nmin0 VDD LPPFET W=1.28U L=0.12U M=1 
X7 nmin0 A VSS VSS LPNFET W=0.76U L=0.12U M=1 
X8 VDD B nmin1 VDD LPPFET W=1.28U L=0.12U M=1 
X9 nmin1 B VSS VSS LPNFET W=0.92U L=0.12U M=1 
.ENDS MX2X8TS 

**** 
*.SUBCKT MX2XLTS Y A B S0 
.SUBCKT MX2XLTS Y A B S0 VSS VDD
X0 net25 nmsel nmin0 VSS LPNFET W=0.2U L=0.12U M=1 
X1 net25 S0 nmin1 VSS LPNFET W=0.2U L=0.12U M=1 
X10 VDD S0 nmsel VDD LPPFET W=0.28U L=0.12U M=1 
X11 nmsel S0 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 net25 S0 nmin0 VDD LPPFET W=0.28U L=0.12U M=1 
X3 net25 nmsel nmin1 VDD LPPFET W=0.28U L=0.12U M=1 
X4 VDD net25 Y VDD LPPFET W=0.42U L=0.12U M=1 
X5 Y net25 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X6 VDD A nmin0 VDD LPPFET W=0.28U L=0.12U M=1 
X7 nmin0 A VSS VSS LPNFET W=0.2U L=0.12U M=1 
X8 VDD B nmin1 VDD LPPFET W=0.28U L=0.12U M=1 
X9 nmin1 B VSS VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS MX2XLTS 

**** 
*.SUBCKT MX3X1TS Y A B C S0 S1 
.SUBCKT MX3X1TS Y A B C S0 S1 VSS VDD
X0 net43 nmsel0 nmin0 VSS LPNFET W=0.56U L=0.12U M=1 
X1 net43 S0 nmin1 VSS LPNFET W=0.56U L=0.12U M=1 
X10 VDD B nmin1 VDD LPPFET W=0.78U L=0.12U M=1 
X11 nmin1 B VSS VSS LPNFET W=0.56U L=0.12U M=1 
X12 VDD C nmin2 VDD LPPFET W=0.5U L=0.12U M=1 
X13 nmin2 C VSS VSS LPNFET W=0.36U L=0.12U M=1 
X14 VDD S0 nmsel0 VDD LPPFET W=0.3U L=0.12U M=1 
X15 nmsel0 S0 VSS VSS LPNFET W=0.22U L=0.12U M=1 
X16 VDD net49 Y VDD LPPFET W=0.64U L=0.12U M=1 
X17 Y net49 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X18 VDD S1 nmsel1 VDD LPPFET W=0.28U L=0.12U M=1 
X19 nmsel1 S1 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 net49 nmsel1 net43 VSS LPNFET W=0.56U L=0.12U M=1 
X3 net49 S1 nmin2 VSS LPNFET W=0.36U L=0.12U M=1 
X4 net43 S0 nmin0 VDD LPPFET W=0.78U L=0.12U M=1 
X5 net43 nmsel0 nmin1 VDD LPPFET W=0.78U L=0.12U M=1 
X6 net49 S1 net43 VDD LPPFET W=0.78U L=0.12U M=1 
X7 net49 nmsel1 nmin2 VDD LPPFET W=0.5U L=0.12U M=1 
X8 VDD A nmin0 VDD LPPFET W=0.78U L=0.12U M=1 
X9 nmin0 A VSS VSS LPNFET W=0.56U L=0.12U M=1 
.ENDS MX3X1TS 

**** 
*.SUBCKT MX3X2TS Y A B C S0 S1 
.SUBCKT MX3X2TS Y A B C S0 S1 VSS VDD
X0 net43 nmsel0 nmin0 VSS LPNFET W=0.86U L=0.12U M=1 
X1 net43 S0 nmin1 VSS LPNFET W=0.86U L=0.12U M=1 
X10 VDD B nmin1 VDD LPPFET W=1.28U L=0.12U M=1 
X11 nmin1 B VSS VSS LPNFET W=0.86U L=0.12U M=1 
X12 VDD C nmin2 VDD LPPFET W=1.02U L=0.12U M=1 
X13 nmin2 C VSS VSS LPNFET W=0.74U L=0.12U M=1 
X14 VDD S0 nmsel0 VDD LPPFET W=0.5U L=0.12U M=1 
X15 nmsel0 S0 VSS VSS LPNFET W=0.36U L=0.12U M=1 
X16 VDD net49 Y VDD LPPFET W=1.28U L=0.12U M=1 
X17 Y net49 VSS VSS LPNFET W=0.86U L=0.12U M=1 
X18 VDD S1 nmsel1 VDD LPPFET W=0.44U L=0.12U M=1 
X19 nmsel1 S1 VSS VSS LPNFET W=0.32U L=0.12U M=1 
X2 net49 nmsel1 net43 VSS LPNFET W=0.86U L=0.12U M=1 
X3 net49 S1 nmin2 VSS LPNFET W=0.74U L=0.12U M=1 
X4 net43 S0 nmin0 VDD LPPFET W=1.28U L=0.12U M=1 
X5 net43 nmsel0 nmin1 VDD LPPFET W=1.28U L=0.12U M=1 
X6 net49 S1 net43 VDD LPPFET W=1.28U L=0.12U M=1 
X7 net49 nmsel1 nmin2 VDD LPPFET W=1.02U L=0.12U M=1 
X8 VDD A nmin0 VDD LPPFET W=1.28U L=0.12U M=1 
X9 nmin0 A VSS VSS LPNFET W=0.86U L=0.12U M=1 
.ENDS MX3X2TS 

**** 
*.SUBCKT MX3X4TS Y A B C S0 S1 
.SUBCKT MX3X4TS Y A B C S0 S1 VSS VDD
X0 net43 nmsel0 nmin0 VSS LPNFET W=0.86U L=0.12U M=1 
X1 net43 S0 nmin1 VSS LPNFET W=0.86U L=0.12U M=1 
X10 VDD B nmin1 VDD LPPFET W=1.28U L=0.12U M=1 
X11 nmin1 B VSS VSS LPNFET W=0.86U L=0.12U M=1 
X12 VDD C nmin2 VDD LPPFET W=1.28U L=0.12U M=1 
X13 nmin2 C VSS VSS LPNFET W=0.92U L=0.12U M=1 
X14 VDD S0 nmsel0 VDD LPPFET W=0.5U L=0.12U M=1 
X15 nmsel0 S0 VSS VSS LPNFET W=0.36U L=0.12U M=1 
X16 VDD net49 Y VDD LPPFET W=2.56U L=0.12U M=1 
X17 Y net49 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X18 VDD S1 nmsel1 VDD LPPFET W=0.46U L=0.12U M=1 
X19 nmsel1 S1 VSS VSS LPNFET W=0.36U L=0.12U M=1 
X2 net49 nmsel1 net43 VSS LPNFET W=0.88U L=0.12U M=1 
X3 net49 S1 nmin2 VSS LPNFET W=0.88U L=0.12U M=1 
X4 net43 S0 nmin0 VDD LPPFET W=1.28U L=0.12U M=1 
X5 net43 nmsel0 nmin1 VDD LPPFET W=1.28U L=0.12U M=1 
X6 net49 S1 net43 VDD LPPFET W=1.28U L=0.12U M=1 
X7 net49 nmsel1 nmin2 VDD LPPFET W=1.28U L=0.12U M=1 
X8 VDD A nmin0 VDD LPPFET W=1.28U L=0.12U M=1 
X9 nmin0 A VSS VSS LPNFET W=0.86U L=0.12U M=1 
.ENDS MX3X4TS 

**** 
*.SUBCKT MX3XLTS Y A B C S0 S1 
.SUBCKT MX3XLTS Y A B C S0 S1 VSS VDD
X0 net43 nmsel0 nmin0 VSS LPNFET W=0.32U L=0.12U M=1 
X1 net43 S0 nmin1 VSS LPNFET W=0.32U L=0.12U M=1 
X10 VDD B nmin1 VDD LPPFET W=0.28U L=0.12U M=1 
X11 nmin1 B VSS VSS LPNFET W=0.2U L=0.12U M=1 
X12 VDD C nmin2 VDD LPPFET W=0.28U L=0.12U M=1 
X13 nmin2 C VSS VSS LPNFET W=0.2U L=0.12U M=1 
X14 VDD S0 nmsel0 VDD LPPFET W=0.28U L=0.12U M=1 
X15 nmsel0 S0 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X16 VDD net49 Y VDD LPPFET W=0.42U L=0.12U M=1 
X17 Y net49 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X18 VDD S1 nmsel1 VDD LPPFET W=0.28U L=0.12U M=1 
X19 nmsel1 S1 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 net49 nmsel1 net43 VSS LPNFET W=0.32U L=0.12U M=1 
X3 net49 S1 nmin2 VSS LPNFET W=0.32U L=0.12U M=1 
X4 net43 S0 nmin0 VDD LPPFET W=0.56U L=0.12U M=1 
X5 net43 nmsel0 nmin1 VDD LPPFET W=0.56U L=0.12U M=1 
X6 net49 S1 net43 VDD LPPFET W=0.56U L=0.12U M=1 
X7 net49 nmsel1 nmin2 VDD LPPFET W=0.56U L=0.12U M=1 
X8 VDD A nmin0 VDD LPPFET W=0.28U L=0.12U M=1 
X9 nmin0 A VSS VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS MX3XLTS 

**** 
*.SUBCKT MX4X1TS Y A B C D S0 S1 
.SUBCKT MX4X1TS Y A B C D S0 S1 VSS VDD
X0 net56 nmsel0 nmin0 VSS LPNFET W=0.54U L=0.12U M=1 
X1 net56 S0 nmin1 VSS LPNFET W=0.54U L=0.12U M=1 
X10 net68 S1 net56 VDD LPPFET W=0.74U L=0.12U M=1 
X11 net68 nmsel1 net62 VDD LPPFET W=0.74U L=0.12U M=1 
X12 VDD A nmin0 VDD LPPFET W=0.78U L=0.12U M=1 
X13 nmin0 A VSS VSS LPNFET W=0.54U L=0.12U M=1 
X14 VDD B nmin1 VDD LPPFET W=0.72U L=0.12U M=1 
X15 nmin1 B VSS VSS LPNFET W=0.54U L=0.12U M=1 
X16 VDD C nmin2 VDD LPPFET W=0.74U L=0.12U M=1 
X17 nmin2 C VSS VSS LPNFET W=0.5U L=0.12U M=1 
X18 VDD D nmin3 VDD LPPFET W=0.74U L=0.12U M=1 
X19 nmin3 D VSS VSS LPNFET W=0.5U L=0.12U M=1 
X2 net62 nmsel0 nmin2 VSS LPNFET W=0.5U L=0.12U M=1 
X20 VDD S0 nmsel0 VDD LPPFET W=0.62U L=0.12U M=1 
X21 nmsel0 S0 VSS VSS LPNFET W=0.44U L=0.12U M=1 
X22 VDD net68 Y VDD LPPFET W=0.64U L=0.12U M=1 
X23 Y net68 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X24 VDD S1 nmsel1 VDD LPPFET W=0.3U L=0.12U M=1 
X25 nmsel1 S1 VSS VSS LPNFET W=0.22U L=0.12U M=1 
X3 net62 S0 nmin3 VSS LPNFET W=0.5U L=0.12U M=1 
X4 net68 nmsel1 net56 VSS LPNFET W=0.5U L=0.12U M=1 
X5 net68 S1 net62 VSS LPNFET W=0.5U L=0.12U M=1 
X6 net56 S0 nmin0 VDD LPPFET W=0.72U L=0.12U M=1 
X7 net56 nmsel0 nmin1 VDD LPPFET W=0.72U L=0.12U M=1 
X8 net62 S0 nmin2 VDD LPPFET W=0.74U L=0.12U M=1 
X9 net62 nmsel0 nmin3 VDD LPPFET W=0.74U L=0.12U M=1 
.ENDS MX4X1TS 

**** 
*.SUBCKT MX4X2TS Y A B C D S0 S1 
.SUBCKT MX4X2TS Y A B C D S0 S1 VSS VDD
X0 net56 nmsel0 nmin0 VSS LPNFET W=0.88U L=0.12U M=1 
X1 net56 S0 nmin1 VSS LPNFET W=0.88U L=0.12U M=1 
X10 net68 S1 net56 VDD LPPFET W=1.24U L=0.12U M=1 
X11 net68 nmsel1 net62 VDD LPPFET W=1.24U L=0.12U M=1 
X12 VDD A nmin0 VDD LPPFET W=1.28U L=0.12U M=1 
X13 nmin0 A VSS VSS LPNFET W=0.88U L=0.12U M=1 
X14 VDD B nmin1 VDD LPPFET W=1.28U L=0.12U M=1 
X15 nmin1 B VSS VSS LPNFET W=0.88U L=0.12U M=1 
X16 VDD C nmin2 VDD LPPFET W=1.24U L=0.12U M=1 
X17 nmin2 C VSS VSS LPNFET W=0.92U L=0.12U M=1 
X18 VDD D nmin3 VDD LPPFET W=1.24U L=0.12U M=1 
X19 nmin3 D VSS VSS LPNFET W=0.92U L=0.12U M=1 
X2 net62 nmsel0 nmin2 VSS LPNFET W=0.92U L=0.12U M=1 
X20 VDD S0 nmsel0 VDD LPPFET W=1.02U L=0.12U M=1 
X21 nmsel0 S0 VSS VSS LPNFET W=0.72U L=0.12U M=1 
X22 VDD net68 Y VDD LPPFET W=1.28U L=0.12U M=1 
X23 Y net68 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X24 VDD S1 nmsel1 VDD LPPFET W=0.5U L=0.12U M=1 
X25 nmsel1 S1 VSS VSS LPNFET W=0.36U L=0.12U M=1 
X3 net62 S0 nmin3 VSS LPNFET W=0.92U L=0.12U M=1 
X4 net68 nmsel1 net56 VSS LPNFET W=0.92U L=0.12U M=1 
X5 net68 S1 net62 VSS LPNFET W=0.92U L=0.12U M=1 
X6 net56 S0 nmin0 VDD LPPFET W=1.28U L=0.12U M=1 
X7 net56 nmsel0 nmin1 VDD LPPFET W=1.28U L=0.12U M=1 
X8 net62 S0 nmin2 VDD LPPFET W=1.24U L=0.12U M=1 
X9 net62 nmsel0 nmin3 VDD LPPFET W=1.24U L=0.12U M=1 
.ENDS MX4X2TS 

**** 
*.SUBCKT MX4X4TS Y A B C D S0 S1 
.SUBCKT MX4X4TS Y A B C D S0 S1 VSS VDD
X0 net56 nmsel0 nmin0 VSS LPNFET W=0.88U L=0.12U M=1 
X1 net56 S0 nmin1 VSS LPNFET W=0.88U L=0.12U M=1 
X10 net68 S1 net56 VDD LPPFET W=1.24U L=0.12U M=1 
X11 net68 nmsel1 net62 VDD LPPFET W=1.24U L=0.12U M=1 
X12 VDD A nmin0 VDD LPPFET W=1.28U L=0.12U M=1 
X13 nmin0 A VSS VSS LPNFET W=0.88U L=0.12U M=1 
X14 VDD B nmin1 VDD LPPFET W=1.28U L=0.12U M=1 
X15 nmin1 B VSS VSS LPNFET W=0.88U L=0.12U M=1 
X16 VDD C nmin2 VDD LPPFET W=1.24U L=0.12U M=1 
X17 nmin2 C VSS VSS LPNFET W=0.92U L=0.12U M=1 
X18 VDD D nmin3 VDD LPPFET W=1.24U L=0.12U M=1 
X19 nmin3 D VSS VSS LPNFET W=0.92U L=0.12U M=1 
X2 net62 nmsel0 nmin2 VSS LPNFET W=0.92U L=0.12U M=1 
X20 VDD S0 nmsel0 VDD LPPFET W=0.98U L=0.12U M=1 
X21 nmsel0 S0 VSS VSS LPNFET W=0.7U L=0.12U M=1 
X22 VDD net68 Y VDD LPPFET W=2.56U L=0.12U M=1 
X23 Y net68 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X24 VDD S1 nmsel1 VDD LPPFET W=0.5U L=0.12U M=1 
X25 nmsel1 S1 VSS VSS LPNFET W=0.36U L=0.12U M=1 
X3 net62 S0 nmin3 VSS LPNFET W=0.92U L=0.12U M=1 
X4 net68 nmsel1 net56 VSS LPNFET W=0.92U L=0.12U M=1 
X5 net68 S1 net62 VSS LPNFET W=0.92U L=0.12U M=1 
X6 net56 S0 nmin0 VDD LPPFET W=1.28U L=0.12U M=1 
X7 net56 nmsel0 nmin1 VDD LPPFET W=1.28U L=0.12U M=1 
X8 net62 S0 nmin2 VDD LPPFET W=1.24U L=0.12U M=1 
X9 net62 nmsel0 nmin3 VDD LPPFET W=1.24U L=0.12U M=1 
.ENDS MX4X4TS 

**** 
*.SUBCKT MX4XLTS Y A B C D S0 S1 
.SUBCKT MX4XLTS Y A B C D S0 S1 VSS VDD
X0 net56 nmsel0 nmin0 VSS LPNFET W=0.2U L=0.12U M=1 
X1 net56 S0 nmin1 VSS LPNFET W=0.2U L=0.12U M=1 
X10 net68 S1 net56 VDD LPPFET W=0.28U L=0.12U M=1 
X11 net68 nmsel1 net62 VDD LPPFET W=0.28U L=0.12U M=1 
X12 VDD A nmin0 VDD LPPFET W=0.28U L=0.12U M=1 
X13 nmin0 A VSS VSS LPNFET W=0.2U L=0.12U M=1 
X14 VDD B nmin1 VDD LPPFET W=0.28U L=0.12U M=1 
X15 nmin1 B VSS VSS LPNFET W=0.18U L=0.12U M=1 
X16 VDD C nmin2 VDD LPPFET W=0.28U L=0.12U M=1 
X17 nmin2 C VSS VSS LPNFET W=0.2U L=0.12U M=1 
X18 VDD D nmin3 VDD LPPFET W=0.28U L=0.12U M=1 
X19 nmin3 D VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 net62 nmsel0 nmin2 VSS LPNFET W=0.2U L=0.12U M=1 
X20 VDD S0 nmsel0 VDD LPPFET W=0.28U L=0.12U M=1 
X21 nmsel0 S0 VSS VSS LPNFET W=0.18U L=0.12U M=1 
X22 VDD net68 Y VDD LPPFET W=0.42U L=0.12U M=1 
X23 Y net68 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X24 VDD S1 nmsel1 VDD LPPFET W=0.28U L=0.12U M=1 
X25 nmsel1 S1 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 net62 S0 nmin3 VSS LPNFET W=0.2U L=0.12U M=1 
X4 net68 nmsel1 net56 VSS LPNFET W=0.2U L=0.12U M=1 
X5 net68 S1 net62 VSS LPNFET W=0.2U L=0.12U M=1 
X6 net56 S0 nmin0 VDD LPPFET W=0.28U L=0.12U M=1 
X7 net56 nmsel0 nmin1 VDD LPPFET W=0.28U L=0.12U M=1 
X8 net62 S0 nmin2 VDD LPPFET W=0.26U L=0.12U M=1 
X9 net62 nmsel0 nmin3 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS MX4XLTS 

**** 
*.SUBCKT MXI2X1TS Y A B S0 
.SUBCKT MXI2X1TS Y A B S0 VSS VDD
X0 Y nmsel nmin0 VSS LPNFET W=0.46U L=0.12U M=1 
X1 Y S0 nmin1 VSS LPNFET W=0.46U L=0.12U M=1 
X2 Y S0 nmin0 VDD LPPFET W=0.64U L=0.12U M=1 
X3 Y nmsel nmin1 VDD LPPFET W=0.64U L=0.12U M=1 
X4 VDD A nmin0 VDD LPPFET W=0.64U L=0.12U M=1 
X5 nmin0 A VSS VSS LPNFET W=0.46U L=0.12U M=1 
X6 VDD B nmin1 VDD LPPFET W=0.64U L=0.12U M=1 
X7 nmin1 B VSS VSS LPNFET W=0.46U L=0.12U M=1 
X8 VDD S0 nmsel VDD LPPFET W=0.28U L=0.12U M=1 
X9 nmsel S0 VSS VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS MXI2X1TS 

**** 
*.SUBCKT MXI2X2TS Y A B S0 
.SUBCKT MXI2X2TS Y A B S0 VSS VDD
X0 Y nmsel nmin0 VSS LPNFET W=0.92U L=0.12U M=1 
X1 Y S0 nmin1 VSS LPNFET W=0.92U L=0.12U M=1 
X2 Y S0 nmin0 VDD LPPFET W=1.2U L=0.12U M=1 
X3 Y nmsel nmin1 VDD LPPFET W=1.2U L=0.12U M=1 
X4 VDD A nmin0 VDD LPPFET W=1.2U L=0.12U M=1 
X5 nmin0 A VSS VSS LPNFET W=0.92U L=0.12U M=1 
X6 VDD B nmin1 VDD LPPFET W=1.16U L=0.12U M=1 
X7 nmin1 B VSS VSS LPNFET W=0.72U L=0.12U M=1 
X8 VDD S0 nmsel VDD LPPFET W=0.5U L=0.12U M=1 
X9 nmsel S0 VSS VSS LPNFET W=0.36U L=0.12U M=1 
.ENDS MXI2X2TS 

**** 
*.SUBCKT MXI2X4TS Y A B S0 
.SUBCKT MXI2X4TS Y A B S0 VSS VDD
X0 Y nmsel nmin0 VSS LPNFET W=1.82U L=0.12U M=1 
X1 Y S0 nmin1 VSS LPNFET W=1.82U L=0.12U M=1 
X2 Y S0 nmin0 VDD LPPFET W=2.44U L=0.12U M=1 
X3 Y nmsel nmin1 VDD LPPFET W=2.44U L=0.12U M=1 
X4 VDD A nmin0 VDD LPPFET W=2.56U L=0.12U M=1 
X5 nmin0 A VSS VSS LPNFET W=1.84U L=0.12U M=1 
X6 VDD B nmin1 VDD LPPFET W=2.56U L=0.12U M=1 
X7 nmin1 B VSS VSS LPNFET W=1.84U L=0.12U M=1 
X8 VDD S0 nmsel VDD LPPFET W=1.02U L=0.12U M=1 
X9 nmsel S0 VSS VSS LPNFET W=0.74U L=0.12U M=1 
.ENDS MXI2X4TS 

**** 
*.SUBCKT MXI2X6TS Y A B S0 
.SUBCKT MXI2X6TS Y A B S0 VSS VDD
X0 hnet20 B VSS VSS LPNFET W=0.46U L=0.12U M=1 
X1 hnet10 B VSS VSS LPNFET W=0.46U L=0.12U M=1 
X10 Y S0 hnet24 VSS LPNFET W=0.46U L=0.12U M=1 
X11 Y S0 hnet18 VSS LPNFET W=0.46U L=0.12U M=1 
X12 hnet23 nmsel Y VDD LPPFET W=0.64U L=0.12U M=1 
X13 hnet21 nmsel Y VDD LPPFET W=0.64U L=0.12U M=1 
X14 hnet25 nmsel Y VDD LPPFET W=0.64U L=0.12U M=1 
X15 hnet12 nmsel Y VDD LPPFET W=0.64U L=0.12U M=1 
X16 hnet14 nmsel Y VDD LPPFET W=0.64U L=0.12U M=1 
X17 hnet9 nmsel Y VDD LPPFET W=0.64U L=0.12U M=1 
X18 VDD B hnet23 VDD LPPFET W=0.64U L=0.12U M=1 
X19 VDD B hnet21 VDD LPPFET W=0.64U L=0.12U M=1 
X2 hnet13 B VSS VSS LPNFET W=0.46U L=0.12U M=1 
X20 VDD B hnet25 VDD LPPFET W=0.64U L=0.12U M=1 
X21 VDD B hnet12 VDD LPPFET W=0.64U L=0.12U M=1 
X22 VDD B hnet14 VDD LPPFET W=0.64U L=0.12U M=1 
X23 VDD B hnet9 VDD LPPFET W=0.64U L=0.12U M=1 
X24 hnet38 A VSS VSS LPNFET W=0.46U L=0.12U M=1 
X25 hnet28 A VSS VSS LPNFET W=0.46U L=0.12U M=1 
X26 hnet31 A VSS VSS LPNFET W=0.46U L=0.12U M=1 
X27 hnet29 A VSS VSS LPNFET W=0.46U L=0.12U M=1 
X28 hnet42 A VSS VSS LPNFET W=0.46U L=0.12U M=1 
X29 hnet36 A VSS VSS LPNFET W=0.46U L=0.12U M=1 
X3 hnet11 B VSS VSS LPNFET W=0.46U L=0.12U M=1 
X30 Y nmsel hnet38 VSS LPNFET W=0.46U L=0.12U M=1 
X31 Y nmsel hnet28 VSS LPNFET W=0.46U L=0.12U M=1 
X32 Y nmsel hnet31 VSS LPNFET W=0.46U L=0.12U M=1 
X33 Y nmsel hnet29 VSS LPNFET W=0.46U L=0.12U M=1 
X34 Y nmsel hnet42 VSS LPNFET W=0.46U L=0.12U M=1 
X35 Y nmsel hnet36 VSS LPNFET W=0.46U L=0.12U M=1 
X36 hnet41 S0 Y VDD LPPFET W=0.64U L=0.12U M=1 
X37 hnet39 S0 Y VDD LPPFET W=0.64U L=0.12U M=1 
X38 hnet43 S0 Y VDD LPPFET W=0.64U L=0.12U M=1 
X39 hnet30 S0 Y VDD LPPFET W=0.64U L=0.12U M=1 
X4 hnet24 B VSS VSS LPNFET W=0.46U L=0.12U M=1 
X40 hnet32 S0 Y VDD LPPFET W=0.64U L=0.12U M=1 
X41 hnet27 S0 Y VDD LPPFET W=0.64U L=0.12U M=1 
X42 VDD A hnet41 VDD LPPFET W=0.64U L=0.12U M=1 
X43 VDD A hnet39 VDD LPPFET W=0.64U L=0.12U M=1 
X44 VDD A hnet43 VDD LPPFET W=0.64U L=0.12U M=1 
X45 VDD A hnet30 VDD LPPFET W=0.64U L=0.12U M=1 
X46 VDD A hnet32 VDD LPPFET W=0.64U L=0.12U M=1 
X47 VDD A hnet27 VDD LPPFET W=0.64U L=0.12U M=1 
X48 VDD S0 nmsel VDD LPPFET W=1.54U L=0.12U M=1 
X49 nmsel S0 VSS VSS LPNFET W=1.1U L=0.12U M=1 
X5 hnet18 B VSS VSS LPNFET W=0.46U L=0.12U M=1 
X6 Y S0 hnet20 VSS LPNFET W=0.46U L=0.12U M=1 
X7 Y S0 hnet10 VSS LPNFET W=0.46U L=0.12U M=1 
X8 Y S0 hnet13 VSS LPNFET W=0.46U L=0.12U M=1 
X9 Y S0 hnet11 VSS LPNFET W=0.46U L=0.12U M=1 
.ENDS MXI2X6TS 

**** 
*.SUBCKT MXI2X8TS Y A B S0 
.SUBCKT MXI2X8TS Y A B S0 VSS VDD
X0 hnet21 B VSS VSS LPNFET W=0.62U L=0.12U M=1 
X1 hnet24 B VSS VSS LPNFET W=0.62U L=0.12U M=1 
X10 Y S0 hnet23 VSS LPNFET W=0.62U L=0.12U M=1 
X11 Y S0 hnet27 VSS LPNFET W=0.62U L=0.12U M=1 
X12 Y S0 hnet17 VSS LPNFET W=0.62U L=0.12U M=1 
X13 Y S0 hnet12 VSS LPNFET W=0.62U L=0.12U M=1 
X14 Y S0 hnet13 VSS LPNFET W=0.62U L=0.12U M=1 
X15 Y S0 hnet11 VSS LPNFET W=0.62U L=0.12U M=1 
X16 hnet9 nmsel Y VDD LPPFET W=0.86U L=0.12U M=1 
X17 hnet22 nmsel Y VDD LPPFET W=0.86U L=0.12U M=1 
X18 VDD B hnet9 VDD LPPFET W=0.86U L=0.12U M=1 
X19 VDD B hnet22 VDD LPPFET W=0.86U L=0.12U M=1 
X2 Y S0 hnet21 VSS LPNFET W=0.62U L=0.12U M=1 
X20 hnet18 nmsel Y VDD LPPFET W=0.86U L=0.12U M=1 
X21 hnet19 nmsel Y VDD LPPFET W=0.86U L=0.12U M=1 
X22 hnet16 nmsel Y VDD LPPFET W=0.86U L=0.12U M=1 
X23 hnet29 nmsel Y VDD LPPFET W=0.86U L=0.12U M=1 
X24 hnet10 nmsel Y VDD LPPFET W=0.86U L=0.12U M=1 
X25 hnet26 nmsel Y VDD LPPFET W=0.86U L=0.12U M=1 
X26 VDD B hnet18 VDD LPPFET W=0.86U L=0.12U M=1 
X27 VDD B hnet19 VDD LPPFET W=0.86U L=0.12U M=1 
X28 VDD B hnet16 VDD LPPFET W=0.86U L=0.12U M=1 
X29 VDD B hnet29 VDD LPPFET W=0.86U L=0.12U M=1 
X3 Y S0 hnet24 VSS LPNFET W=0.62U L=0.12U M=1 
X30 VDD B hnet10 VDD LPPFET W=0.86U L=0.12U M=1 
X31 VDD B hnet26 VDD LPPFET W=0.86U L=0.12U M=1 
X32 hnet43 A VSS VSS LPNFET W=0.62U L=0.12U M=1 
X33 hnet46 A VSS VSS LPNFET W=0.62U L=0.12U M=1 
X34 Y nmsel hnet43 VSS LPNFET W=0.62U L=0.12U M=1 
X35 Y nmsel hnet46 VSS LPNFET W=0.62U L=0.12U M=1 
X36 hnet45 A VSS VSS LPNFET W=0.62U L=0.12U M=1 
X37 hnet49 A VSS VSS LPNFET W=0.62U L=0.12U M=1 
X38 hnet39 A VSS VSS LPNFET W=0.62U L=0.12U M=1 
X39 hnet34 A VSS VSS LPNFET W=0.62U L=0.12U M=1 
X4 hnet23 B VSS VSS LPNFET W=0.62U L=0.12U M=1 
X40 hnet35 A VSS VSS LPNFET W=0.62U L=0.12U M=1 
X41 hnet33 A VSS VSS LPNFET W=0.62U L=0.12U M=1 
X42 Y nmsel hnet45 VSS LPNFET W=0.62U L=0.12U M=1 
X43 Y nmsel hnet49 VSS LPNFET W=0.62U L=0.12U M=1 
X44 Y nmsel hnet39 VSS LPNFET W=0.62U L=0.12U M=1 
X45 Y nmsel hnet34 VSS LPNFET W=0.62U L=0.12U M=1 
X46 Y nmsel hnet35 VSS LPNFET W=0.62U L=0.12U M=1 
X47 Y nmsel hnet33 VSS LPNFET W=0.62U L=0.12U M=1 
X48 hnet31 S0 Y VDD LPPFET W=0.86U L=0.12U M=1 
X49 hnet44 S0 Y VDD LPPFET W=0.86U L=0.12U M=1 
X5 hnet27 B VSS VSS LPNFET W=0.62U L=0.12U M=1 
X50 VDD A hnet31 VDD LPPFET W=0.86U L=0.12U M=1 
X51 VDD A hnet44 VDD LPPFET W=0.86U L=0.12U M=1 
X52 hnet40 S0 Y VDD LPPFET W=0.86U L=0.12U M=1 
X53 hnet41 S0 Y VDD LPPFET W=0.86U L=0.12U M=1 
X54 hnet38 S0 Y VDD LPPFET W=0.86U L=0.12U M=1 
X55 hnet51 S0 Y VDD LPPFET W=0.86U L=0.12U M=1 
X56 hnet32 S0 Y VDD LPPFET W=0.86U L=0.12U M=1 
X57 hnet48 S0 Y VDD LPPFET W=0.86U L=0.12U M=1 
X58 VDD A hnet40 VDD LPPFET W=0.86U L=0.12U M=1 
X59 VDD A hnet41 VDD LPPFET W=0.86U L=0.12U M=1 
X6 hnet17 B VSS VSS LPNFET W=0.62U L=0.12U M=1 
X60 VDD A hnet38 VDD LPPFET W=0.86U L=0.12U M=1 
X61 VDD A hnet51 VDD LPPFET W=0.86U L=0.12U M=1 
X62 VDD A hnet32 VDD LPPFET W=0.86U L=0.12U M=1 
X63 VDD A hnet48 VDD LPPFET W=0.86U L=0.12U M=1 
X64 VDD S0 nmsel VDD LPPFET W=2.06U L=0.12U M=1 
X65 nmsel S0 VSS VSS LPNFET W=1.48U L=0.12U M=1 
X7 hnet12 B VSS VSS LPNFET W=0.62U L=0.12U M=1 
X8 hnet13 B VSS VSS LPNFET W=0.62U L=0.12U M=1 
X9 hnet11 B VSS VSS LPNFET W=0.62U L=0.12U M=1 
.ENDS MXI2X8TS 

**** 
*.SUBCKT MXI2XLTS Y A B S0 
.SUBCKT MXI2XLTS Y A B S0 VSS VDD
X0 Y nmsel nmin0 VSS LPNFET W=0.2U L=0.12U M=1 
X1 Y S0 nmin1 VSS LPNFET W=0.2U L=0.12U M=1 
X2 Y S0 nmin0 VDD LPPFET W=0.28U L=0.12U M=1 
X3 Y nmsel nmin1 VDD LPPFET W=0.28U L=0.12U M=1 
X4 VDD A nmin0 VDD LPPFET W=0.42U L=0.12U M=1 
X5 nmin0 A VSS VSS LPNFET W=0.24U L=0.12U M=1 
X6 VDD B nmin1 VDD LPPFET W=0.38U L=0.12U M=1 
X7 nmin1 B VSS VSS LPNFET W=0.18U L=0.12U M=1 
X8 VDD S0 nmsel VDD LPPFET W=0.28U L=0.12U M=1 
X9 nmsel S0 VSS VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS MXI2XLTS 

**** 
*.SUBCKT MXI3X1TS Y A B C S0 S1 
.SUBCKT MXI3X1TS Y A B C S0 S1 VSS VDD
X0 net46 nmsel0 nmin0 VSS LPNFET W=0.28U L=0.12U M=1 
X1 net46 S0 nmin1 VSS LPNFET W=0.26U L=0.12U M=1 
X10 VDD B nmin1 VDD LPPFET W=0.38U L=0.12U M=1 
X11 nmin1 B VSS VSS LPNFET W=0.28U L=0.12U M=1 
X12 VDD C nmin2 VDD LPPFET W=0.28U L=0.12U M=1 
X13 nmin2 C VSS VSS LPNFET W=0.2U L=0.12U M=1 
X14 VDD net46 net74 VDD LPPFET W=0.5U L=0.12U M=1 
X15 net74 net46 VSS VSS LPNFET W=0.36U L=0.12U M=1 
X16 VDD nmin2 net76 VDD LPPFET W=0.5U L=0.12U M=1 
X17 net76 nmin2 VSS VSS LPNFET W=0.36U L=0.12U M=1 
X18 VDD S0 nmsel0 VDD LPPFET W=0.28U L=0.12U M=1 
X19 nmsel0 S0 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 net52 nmsel1 net74 VSS LPNFET W=0.36U L=0.12U M=1 
X20 VDD net52 Y VDD LPPFET W=0.62U L=0.12U M=1 
X21 Y net52 VSS VSS LPNFET W=0.42U L=0.12U M=1 
X22 VDD S1 nmsel1 VDD LPPFET W=0.28U L=0.12U M=1 
X23 nmsel1 S1 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 net52 S1 net76 VSS LPNFET W=0.36U L=0.12U M=1 
X4 net46 S0 nmin0 VDD LPPFET W=0.38U L=0.12U M=1 
X5 net46 nmsel0 nmin1 VDD LPPFET W=0.38U L=0.12U M=1 
X6 net52 S1 net74 VDD LPPFET W=0.5U L=0.12U M=1 
X7 net52 nmsel1 net76 VDD LPPFET W=0.5U L=0.12U M=1 
X8 VDD A nmin0 VDD LPPFET W=0.38U L=0.12U M=1 
X9 nmin0 A VSS VSS LPNFET W=0.28U L=0.12U M=1 
.ENDS MXI3X1TS 

**** 
*.SUBCKT MXI3X2TS Y A B C S0 S1 
.SUBCKT MXI3X2TS Y A B C S0 S1 VSS VDD
X0 net46 nmsel0 nmin0 VSS LPNFET W=0.58U L=0.12U M=1 
X1 net46 S0 nmin1 VSS LPNFET W=0.56U L=0.12U M=1 
X10 VDD B nmin1 VDD LPPFET W=0.78U L=0.12U M=1 
X11 nmin1 B VSS VSS LPNFET W=0.56U L=0.12U M=1 
X12 VDD C nmin2 VDD LPPFET W=0.42U L=0.12U M=1 
X13 nmin2 C VSS VSS LPNFET W=0.3U L=0.12U M=1 
X14 VDD net46 net74 VDD LPPFET W=0.92U L=0.12U M=1 
X15 net74 net46 VSS VSS LPNFET W=0.62U L=0.12U M=1 
X16 VDD nmin2 net76 VDD LPPFET W=0.98U L=0.12U M=1 
X17 net76 nmin2 VSS VSS LPNFET W=0.72U L=0.12U M=1 
X18 VDD S0 nmsel0 VDD LPPFET W=0.34U L=0.12U M=1 
X19 nmsel0 S0 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X2 net52 nmsel1 net74 VSS LPNFET W=0.62U L=0.12U M=1 
X20 VDD net52 Y VDD LPPFET W=1.24U L=0.12U M=1 
X21 Y net52 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X22 VDD S1 nmsel1 VDD LPPFET W=0.42U L=0.12U M=1 
X23 nmsel1 S1 VSS VSS LPNFET W=0.3U L=0.12U M=1 
X3 net52 S1 net76 VSS LPNFET W=0.72U L=0.12U M=1 
X4 net46 S0 nmin0 VDD LPPFET W=0.78U L=0.12U M=1 
X5 net46 nmsel0 nmin1 VDD LPPFET W=0.78U L=0.12U M=1 
X6 net52 S1 net74 VDD LPPFET W=1.02U L=0.12U M=1 
X7 net52 nmsel1 net76 VDD LPPFET W=0.98U L=0.12U M=1 
X8 VDD A nmin0 VDD LPPFET W=0.78U L=0.12U M=1 
X9 nmin0 A VSS VSS LPNFET W=0.58U L=0.12U M=1 
.ENDS MXI3X2TS 

**** 
*.SUBCKT MXI3X4TS Y A B C S0 S1 
.SUBCKT MXI3X4TS Y A B C S0 S1 VSS VDD
X0 net46 nmsel0 nmin0 VSS LPNFET W=0.72U L=0.12U M=1 
X1 net46 S0 nmin1 VSS LPNFET W=0.74U L=0.12U M=1 
X10 VDD B nmin1 VDD LPPFET W=0.98U L=0.12U M=1 
X11 nmin1 B VSS VSS LPNFET W=0.6U L=0.12U M=1 
X12 VDD C nmin2 VDD LPPFET W=0.5U L=0.12U M=1 
X13 nmin2 C VSS VSS LPNFET W=0.36U L=0.12U M=1 
X14 VDD net46 net74 VDD LPPFET W=1.28U L=0.12U M=1 
X15 net74 net46 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X16 VDD nmin2 net76 VDD LPPFET W=1.16U L=0.12U M=1 
X17 net76 nmin2 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X18 VDD S0 nmsel0 VDD LPPFET W=0.42U L=0.12U M=1 
X19 nmsel0 S0 VSS VSS LPNFET W=0.3U L=0.12U M=1 
X2 net52 nmsel1 net74 VSS LPNFET W=0.72U L=0.12U M=1 
X20 VDD net52 Y VDD LPPFET W=2.56U L=0.12U M=1 
X21 Y net52 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X22 VDD S1 nmsel1 VDD LPPFET W=0.5U L=0.12U M=1 
X23 nmsel1 S1 VSS VSS LPNFET W=0.36U L=0.12U M=1 
X3 net52 S1 net76 VSS LPNFET W=0.92U L=0.12U M=1 
X4 net46 S0 nmin0 VDD LPPFET W=1.02U L=0.12U M=1 
X5 net46 nmsel0 nmin1 VDD LPPFET W=0.98U L=0.12U M=1 
X6 net52 S1 net74 VDD LPPFET W=1.16U L=0.12U M=1 
X7 net52 nmsel1 net76 VDD LPPFET W=1.16U L=0.12U M=1 
X8 VDD A nmin0 VDD LPPFET W=1.02U L=0.12U M=1 
X9 nmin0 A VSS VSS LPNFET W=0.72U L=0.12U M=1 
.ENDS MXI3X4TS 

**** 
*.SUBCKT MXI3XLTS Y A B C S0 S1 
.SUBCKT MXI3XLTS Y A B C S0 S1 VSS VDD
X0 net46 nmsel0 nmin0 VSS LPNFET W=0.32U L=0.12U M=1 
X1 net46 S0 nmin1 VSS LPNFET W=0.32U L=0.12U M=1 
X10 VDD B nmin1 VDD LPPFET W=0.28U L=0.12U M=1 
X11 nmin1 B VSS VSS LPNFET W=0.2U L=0.12U M=1 
X12 VDD C nmin2 VDD LPPFET W=0.28U L=0.12U M=1 
X13 nmin2 C VSS VSS LPNFET W=0.2U L=0.12U M=1 
X14 VDD net46 net74 VDD LPPFET W=0.28U L=0.12U M=1 
X15 net74 net46 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X16 VDD nmin2 net76 VDD LPPFET W=0.28U L=0.12U M=1 
X17 net76 nmin2 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X18 VDD S0 nmsel0 VDD LPPFET W=0.28U L=0.12U M=1 
X19 nmsel0 S0 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 net52 nmsel1 net74 VSS LPNFET W=0.32U L=0.12U M=1 
X20 VDD net52 Y VDD LPPFET W=0.42U L=0.12U M=1 
X21 Y net52 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X22 VDD S1 nmsel1 VDD LPPFET W=0.28U L=0.12U M=1 
X23 nmsel1 S1 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 net52 S1 net76 VSS LPNFET W=0.32U L=0.12U M=1 
X4 net46 S0 nmin0 VDD LPPFET W=0.56U L=0.12U M=1 
X5 net46 nmsel0 nmin1 VDD LPPFET W=0.56U L=0.12U M=1 
X6 net52 S1 net74 VDD LPPFET W=0.56U L=0.12U M=1 
X7 net52 nmsel1 net76 VDD LPPFET W=0.56U L=0.12U M=1 
X8 VDD A nmin0 VDD LPPFET W=0.28U L=0.12U M=1 
X9 nmin0 A VSS VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS MXI3XLTS 

**** 
*.SUBCKT MXI4X1TS Y A B C D S0 S1 
.SUBCKT MXI4X1TS Y A B C D S0 S1 VSS VDD
X0 net58 nmsel0 nmin0 VSS LPNFET W=0.28U L=0.12U M=1 
X1 net58 S0 nmin1 VSS LPNFET W=0.28U L=0.12U M=1 
X10 net70 S1 net100 VDD LPPFET W=0.5U L=0.12U M=1 
X11 net70 nmsel1 net102 VDD LPPFET W=0.5U L=0.12U M=1 
X12 VDD A nmin0 VDD LPPFET W=0.38U L=0.12U M=1 
X13 nmin0 A VSS VSS LPNFET W=0.28U L=0.12U M=1 
X14 VDD B nmin1 VDD LPPFET W=0.38U L=0.12U M=1 
X15 nmin1 B VSS VSS LPNFET W=0.28U L=0.12U M=1 
X16 VDD C nmin2 VDD LPPFET W=0.38U L=0.12U M=1 
X17 nmin2 C VSS VSS LPNFET W=0.28U L=0.12U M=1 
X18 VDD D nmin3 VDD LPPFET W=0.38U L=0.12U M=1 
X19 nmin3 D VSS VSS LPNFET W=0.28U L=0.12U M=1 
X2 net64 nmsel0 nmin2 VSS LPNFET W=0.28U L=0.12U M=1 
X20 VDD net58 net100 VDD LPPFET W=0.5U L=0.12U M=1 
X21 net100 net58 VSS VSS LPNFET W=0.36U L=0.12U M=1 
X22 VDD net64 net102 VDD LPPFET W=0.5U L=0.12U M=1 
X23 net102 net64 VSS VSS LPNFET W=0.36U L=0.12U M=1 
X24 VDD S0 nmsel0 VDD LPPFET W=0.3U L=0.12U M=1 
X25 nmsel0 S0 VSS VSS LPNFET W=0.22U L=0.12U M=1 
X26 VDD net70 Y VDD LPPFET W=0.64U L=0.12U M=1 
X27 Y net70 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X28 VDD S1 nmsel1 VDD LPPFET W=0.28U L=0.12U M=1 
X29 nmsel1 S1 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 net64 S0 nmin3 VSS LPNFET W=0.28U L=0.12U M=1 
X4 net70 nmsel1 net100 VSS LPNFET W=0.36U L=0.12U M=1 
X5 net70 S1 net102 VSS LPNFET W=0.36U L=0.12U M=1 
X6 net58 S0 nmin0 VDD LPPFET W=0.38U L=0.12U M=1 
X7 net58 nmsel0 nmin1 VDD LPPFET W=0.38U L=0.12U M=1 
X8 net64 S0 nmin2 VDD LPPFET W=0.38U L=0.12U M=1 
X9 net64 nmsel0 nmin3 VDD LPPFET W=0.38U L=0.12U M=1 
.ENDS MXI4X1TS 

**** 
*.SUBCKT MXI4X2TS Y A B C D S0 S1 
.SUBCKT MXI4X2TS Y A B C D S0 S1 VSS VDD
X0 net58 nmsel0 nmin0 VSS LPNFET W=0.58U L=0.12U M=1 
X1 net58 S0 nmin1 VSS LPNFET W=0.58U L=0.12U M=1 
X10 net70 S1 net100 VDD LPPFET W=0.92U L=0.12U M=1 
X11 net70 nmsel1 net102 VDD LPPFET W=1.02U L=0.12U M=1 
X12 VDD A nmin0 VDD LPPFET W=0.8U L=0.12U M=1 
X13 nmin0 A VSS VSS LPNFET W=0.58U L=0.12U M=1 
X14 VDD B nmin1 VDD LPPFET W=0.8U L=0.12U M=1 
X15 nmin1 B VSS VSS LPNFET W=0.58U L=0.12U M=1 
X16 VDD C nmin2 VDD LPPFET W=0.76U L=0.12U M=1 
X17 nmin2 C VSS VSS LPNFET W=0.56U L=0.12U M=1 
X18 VDD D nmin3 VDD LPPFET W=0.76U L=0.12U M=1 
X19 nmin3 D VSS VSS LPNFET W=0.54U L=0.12U M=1 
X2 net64 nmsel0 nmin2 VSS LPNFET W=0.58U L=0.12U M=1 
X20 VDD net58 net100 VDD LPPFET W=1.02U L=0.12U M=1 
X21 net100 net58 VSS VSS LPNFET W=0.74U L=0.12U M=1 
X22 VDD net64 net102 VDD LPPFET W=1.02U L=0.12U M=1 
X23 net102 net64 VSS VSS LPNFET W=0.72U L=0.12U M=1 
X24 VDD S0 nmsel0 VDD LPPFET W=0.64U L=0.12U M=1 
X25 nmsel0 S0 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X26 VDD net70 Y VDD LPPFET W=1.28U L=0.12U M=1 
X27 Y net70 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X28 VDD S1 nmsel1 VDD LPPFET W=0.42U L=0.12U M=1 
X29 nmsel1 S1 VSS VSS LPNFET W=0.3U L=0.12U M=1 
X3 net64 S0 nmin3 VSS LPNFET W=0.58U L=0.12U M=1 
X4 net70 nmsel1 net100 VSS LPNFET W=0.68U L=0.12U M=1 
X5 net70 S1 net102 VSS LPNFET W=0.72U L=0.12U M=1 
X6 net58 S0 nmin0 VDD LPPFET W=0.8U L=0.12U M=1 
X7 net58 nmsel0 nmin1 VDD LPPFET W=0.8U L=0.12U M=1 
X8 net64 S0 nmin2 VDD LPPFET W=0.76U L=0.12U M=1 
X9 net64 nmsel0 nmin3 VDD LPPFET W=0.76U L=0.12U M=1 
.ENDS MXI4X2TS 

**** 
*.SUBCKT MXI4X4TS Y A B C D S0 S1 
.SUBCKT MXI4X4TS Y A B C D S0 S1 VSS VDD
X0 net58 nmsel0 nmin0 VSS LPNFET W=0.68U L=0.12U M=1 
X1 net58 S0 nmin1 VSS LPNFET W=0.66U L=0.12U M=1 
X10 net70 S1 net100 VDD LPPFET W=1.16U L=0.12U M=1 
X11 net70 nmsel1 net102 VDD LPPFET W=1.18U L=0.12U M=1 
X12 VDD A nmin0 VDD LPPFET W=1.02U L=0.12U M=1 
X13 nmin0 A VSS VSS LPNFET W=0.68U L=0.12U M=1 
X14 VDD B nmin1 VDD LPPFET W=0.96U L=0.12U M=1 
X15 nmin1 B VSS VSS LPNFET W=0.62U L=0.12U M=1 
X16 VDD C nmin2 VDD LPPFET W=1U L=0.12U M=1 
X17 nmin2 C VSS VSS LPNFET W=0.74U L=0.12U M=1 
X18 VDD D nmin3 VDD LPPFET W=0.96U L=0.12U M=1 
X19 nmin3 D VSS VSS LPNFET W=0.62U L=0.12U M=1 
X2 net64 nmsel0 nmin2 VSS LPNFET W=0.74U L=0.12U M=1 
X20 VDD net58 net100 VDD LPPFET W=1.28U L=0.12U M=1 
X21 net100 net58 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X22 VDD net64 net102 VDD LPPFET W=1.18U L=0.12U M=1 
X23 net102 net64 VSS VSS LPNFET W=0.84U L=0.12U M=1 
X24 VDD S0 nmsel0 VDD LPPFET W=0.8U L=0.12U M=1 
X25 nmsel0 S0 VSS VSS LPNFET W=0.58U L=0.12U M=1 
X26 VDD net70 Y VDD LPPFET W=2.56U L=0.12U M=1 
X27 Y net70 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X28 VDD S1 nmsel1 VDD LPPFET W=0.5U L=0.12U M=1 
X29 nmsel1 S1 VSS VSS LPNFET W=0.36U L=0.12U M=1 
X3 net64 S0 nmin3 VSS LPNFET W=0.74U L=0.12U M=1 
X4 net70 nmsel1 net100 VSS LPNFET W=0.72U L=0.12U M=1 
X5 net70 S1 net102 VSS LPNFET W=0.92U L=0.12U M=1 
X6 net58 S0 nmin0 VDD LPPFET W=1.02U L=0.12U M=1 
X7 net58 nmsel0 nmin1 VDD LPPFET W=0.96U L=0.12U M=1 
X8 net64 S0 nmin2 VDD LPPFET W=1U L=0.12U M=1 
X9 net64 nmsel0 nmin3 VDD LPPFET W=0.96U L=0.12U M=1 
.ENDS MXI4X4TS 

**** 
*.SUBCKT MXI4XLTS Y A B C D S0 S1 
.SUBCKT MXI4XLTS Y A B C D S0 S1 VSS VDD
X0 net58 nmsel0 nmin0 VSS LPNFET W=0.2U L=0.12U M=1 
X1 net58 S0 nmin1 VSS LPNFET W=0.2U L=0.12U M=1 
X10 net70 S1 net100 VDD LPPFET W=0.28U L=0.12U M=1 
X11 net70 nmsel1 net102 VDD LPPFET W=0.28U L=0.12U M=1 
X12 VDD A nmin0 VDD LPPFET W=0.28U L=0.12U M=1 
X13 nmin0 A VSS VSS LPNFET W=0.2U L=0.12U M=1 
X14 VDD B nmin1 VDD LPPFET W=0.28U L=0.12U M=1 
X15 nmin1 B VSS VSS LPNFET W=0.2U L=0.12U M=1 
X16 VDD C nmin2 VDD LPPFET W=0.28U L=0.12U M=1 
X17 nmin2 C VSS VSS LPNFET W=0.2U L=0.12U M=1 
X18 VDD D nmin3 VDD LPPFET W=0.28U L=0.12U M=1 
X19 nmin3 D VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 net64 nmsel0 nmin2 VSS LPNFET W=0.2U L=0.12U M=1 
X20 VDD net58 net100 VDD LPPFET W=0.28U L=0.12U M=1 
X21 net100 net58 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X22 VDD net64 net102 VDD LPPFET W=0.28U L=0.12U M=1 
X23 net102 net64 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X24 VDD S0 nmsel0 VDD LPPFET W=0.28U L=0.12U M=1 
X25 nmsel0 S0 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X26 VDD net70 Y VDD LPPFET W=0.42U L=0.12U M=1 
X27 Y net70 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X28 VDD S1 nmsel1 VDD LPPFET W=0.28U L=0.12U M=1 
X29 nmsel1 S1 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 net64 S0 nmin3 VSS LPNFET W=0.2U L=0.12U M=1 
X4 net70 nmsel1 net100 VSS LPNFET W=0.2U L=0.12U M=1 
X5 net70 S1 net102 VSS LPNFET W=0.2U L=0.12U M=1 
X6 net58 S0 nmin0 VDD LPPFET W=0.28U L=0.12U M=1 
X7 net58 nmsel0 nmin1 VDD LPPFET W=0.28U L=0.12U M=1 
X8 net64 S0 nmin2 VDD LPPFET W=0.28U L=0.12U M=1 
X9 net64 nmsel0 nmin3 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS MXI4XLTS 

**** 
*.SUBCKT NAND2BX1TS Y AN B 
.SUBCKT NAND2BX1TS Y AN B VSS VDD
X0 VDD AN nmin1 VDD LPPFET W=0.28U L=0.12U M=1 
X1 nmin1 AN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 hnet14 B VSS VSS LPNFET W=0.6U L=0.12U M=1 
X3 Y nmin1 hnet14 VSS LPNFET W=0.6U L=0.12U M=1 
X4 VDD B Y VDD LPPFET W=0.64U L=0.12U M=1 
X5 VDD nmin1 Y VDD LPPFET W=0.64U L=0.12U M=1 
.ENDS NAND2BX1TS 

**** 
*.SUBCKT NAND2BX2TS Y AN B 
.SUBCKT NAND2BX2TS Y AN B VSS VDD
X0 VDD AN nmin1 VDD LPPFET W=0.58U L=0.12U M=1 
X1 nmin1 AN VSS VSS LPNFET W=0.42U L=0.12U M=1 
X2 hnet15 B VSS VSS LPNFET W=0.6U L=0.12U M=1 
X3 Y nmin1 hnet15 VSS LPNFET W=0.6U L=0.12U M=1 
X4 hnet11 B VSS VSS LPNFET W=0.6U L=0.12U M=1 
X5 Y nmin1 hnet11 VSS LPNFET W=0.6U L=0.12U M=1 
X6 VDD B Y VDD LPPFET W=1.26U L=0.12U M=1 
X7 VDD nmin1 Y VDD LPPFET W=1.26U L=0.12U M=1 
.ENDS NAND2BX2TS 

**** 
*.SUBCKT NAND2BX4TS Y AN B 
.SUBCKT NAND2BX4TS Y AN B VSS VDD
X0 VDD AN nmin1 VDD LPPFET W=1.16U L=0.12U M=1 
X1 nmin1 AN VSS VSS LPNFET W=0.84U L=0.12U M=1 
X2 hnet11 B VSS VSS LPNFET W=0.82U L=0.12U M=1 
X3 Y nmin1 hnet11 VSS LPNFET W=0.82U L=0.12U M=1 
X4 hnet12 B VSS VSS LPNFET W=0.82U L=0.12U M=1 
X5 Y nmin1 hnet12 VSS LPNFET W=0.82U L=0.12U M=1 
X6 hnet14 B VSS VSS LPNFET W=0.82U L=0.12U M=1 
X7 Y nmin1 hnet14 VSS LPNFET W=0.82U L=0.12U M=1 
X8 VDD B Y VDD LPPFET W=2.44U L=0.12U M=1 
X9 VDD nmin1 Y VDD LPPFET W=2.44U L=0.12U M=1 
.ENDS NAND2BX4TS 

**** 
*.SUBCKT NAND2BXLTS Y AN B 
.SUBCKT NAND2BXLTS Y AN B VSS VDD
X0 VDD AN nmin1 VDD LPPFET W=0.28U L=0.12U M=1 
X1 nmin1 AN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 hnet14 B VSS VSS LPNFET W=0.4U L=0.12U M=1 
X3 Y nmin1 hnet14 VSS LPNFET W=0.4U L=0.12U M=1 
X4 VDD B Y VDD LPPFET W=0.42U L=0.12U M=1 
X5 VDD nmin1 Y VDD LPPFET W=0.42U L=0.12U M=1 
.ENDS NAND2BXLTS 

**** 
*.SUBCKT NAND2X1TS Y A B 
.SUBCKT NAND2X1TS Y A B VSS VDD
X0 hnet11 B VSS VSS LPNFET W=0.6U L=0.12U M=1 
X1 Y A hnet11 VSS LPNFET W=0.6U L=0.12U M=1 
X2 VDD B Y VDD LPPFET W=0.64U L=0.12U M=1 
X3 VDD A Y VDD LPPFET W=0.64U L=0.12U M=1 
.ENDS NAND2X1TS 

**** 
*.SUBCKT NAND2X2TS Y A B 
.SUBCKT NAND2X2TS Y A B VSS VDD
X0 hnet12 B VSS VSS LPNFET W=0.6U L=0.12U M=1 
X1 Y A hnet12 VSS LPNFET W=0.6U L=0.12U M=1 
X2 hnet6 B VSS VSS LPNFET W=0.6U L=0.12U M=1 
X3 Y A hnet6 VSS LPNFET W=0.6U L=0.12U M=1 
X4 VDD B Y VDD LPPFET W=1.26U L=0.12U M=1 
X5 VDD A Y VDD LPPFET W=1.26U L=0.12U M=1 
.ENDS NAND2X2TS 

**** 
*.SUBCKT NAND2X4TS Y A B 
.SUBCKT NAND2X4TS Y A B VSS VDD
X0 net12 B VSS VSS LPNFET W=0.72U L=0.12U M=1 
X1 Y A net12 VSS LPNFET W=0.72U L=0.12U M=1 
X2 net20 B VSS VSS LPNFET W=0.82U L=0.12U M=1 
X3 Y A net20 VSS LPNFET W=0.82U L=0.12U M=1 
X4 net26 B VSS VSS LPNFET W=0.82U L=0.12U M=1 
X5 Y A net26 VSS LPNFET W=0.82U L=0.12U M=1 
X6 VDD B Y VDD LPPFET W=2.58U L=0.12U M=1 
X7 VDD A Y VDD LPPFET W=2.58U L=0.12U M=1 
.ENDS NAND2X4TS 

**** 
*.SUBCKT NAND2X6TS Y A B 
.SUBCKT NAND2X6TS Y A B VSS VDD
X0 hnet14 B VSS VSS LPNFET W=0.86U L=0.12U M=1 
X1 Y A hnet14 VSS LPNFET W=0.86U L=0.12U M=1 
X2 hnet7 B VSS VSS LPNFET W=0.86U L=0.12U M=1 
X3 Y A hnet7 VSS LPNFET W=0.86U L=0.12U M=1 
X4 hnet9 B VSS VSS LPNFET W=0.86U L=0.12U M=1 
X5 Y A hnet9 VSS LPNFET W=0.86U L=0.12U M=1 
X6 hnet13 B VSS VSS LPNFET W=0.86U L=0.12U M=1 
X7 Y A hnet13 VSS LPNFET W=0.86U L=0.12U M=1 
X8 VDD B Y VDD LPPFET W=3.84U L=0.12U M=1 
X9 VDD A Y VDD LPPFET W=3.84U L=0.12U M=1 
.ENDS NAND2X6TS 

**** 
*.SUBCKT NAND2X8TS Y A B 
.SUBCKT NAND2X8TS Y A B VSS VDD
X0 hnet15 B VSS VSS LPNFET W=0.88U L=0.12U M=1 
X1 Y A hnet15 VSS LPNFET W=0.88U L=0.12U M=1 
X10 VDD B Y VDD LPPFET W=4.84U L=0.12U M=1 
X11 VDD A Y VDD LPPFET W=4.84U L=0.12U M=1 
X2 hnet7 B VSS VSS LPNFET W=0.88U L=0.12U M=1 
X3 Y A hnet7 VSS LPNFET W=0.88U L=0.12U M=1 
X4 hnet10 B VSS VSS LPNFET W=0.88U L=0.12U M=1 
X5 Y A hnet10 VSS LPNFET W=0.88U L=0.12U M=1 
X6 hnet14 B VSS VSS LPNFET W=0.88U L=0.12U M=1 
X7 Y A hnet14 VSS LPNFET W=0.88U L=0.12U M=1 
X8 hnet6 B VSS VSS LPNFET W=0.88U L=0.12U M=1 
X9 Y A hnet6 VSS LPNFET W=0.88U L=0.12U M=1 
.ENDS NAND2X8TS 

**** 
*.SUBCKT NAND2XLTS Y A B 
.SUBCKT NAND2XLTS Y A B VSS VDD
X0 hnet11 B VSS VSS LPNFET W=0.4U L=0.12U M=1 
X1 Y A hnet11 VSS LPNFET W=0.4U L=0.12U M=1 
X2 VDD B Y VDD LPPFET W=0.42U L=0.12U M=1 
X3 VDD A Y VDD LPPFET W=0.42U L=0.12U M=1 
.ENDS NAND2XLTS 

**** 
*.SUBCKT NAND3BX1TS Y AN B C 
.SUBCKT NAND3BX1TS Y AN B C VSS VDD
X0 VDD AN nmin1 VDD LPPFET W=0.3U L=0.12U M=1 
X1 nmin1 AN VSS VSS LPNFET W=0.22U L=0.12U M=1 
X2 hnet17 C VSS VSS LPNFET W=0.72U L=0.12U M=1 
X3 hnet12 B hnet17 VSS LPNFET W=0.72U L=0.12U M=1 
X4 Y nmin1 hnet12 VSS LPNFET W=0.72U L=0.12U M=1 
X5 VDD C Y VDD LPPFET W=0.64U L=0.12U M=1 
X6 VDD B Y VDD LPPFET W=0.64U L=0.12U M=1 
X7 VDD nmin1 Y VDD LPPFET W=0.64U L=0.12U M=1 
.ENDS NAND3BX1TS 

**** 
*.SUBCKT NAND3BX2TS Y AN B C 
.SUBCKT NAND3BX2TS Y AN B C VSS VDD
X0 VDD AN nmin1 VDD LPPFET W=0.64U L=0.12U M=1 
X1 nmin1 AN VSS VSS LPNFET W=0.46U L=0.12U M=1 
X10 VDD nmin1 Y VDD LPPFET W=1.14U L=0.12U M=1 
X2 hnet18 C VSS VSS LPNFET W=0.64U L=0.12U M=1 
X3 hnet12 B hnet18 VSS LPNFET W=0.64U L=0.12U M=1 
X4 Y nmin1 hnet12 VSS LPNFET W=0.64U L=0.12U M=1 
X5 hnet19 C VSS VSS LPNFET W=0.64U L=0.12U M=1 
X6 hnet14 B hnet19 VSS LPNFET W=0.64U L=0.12U M=1 
X7 Y nmin1 hnet14 VSS LPNFET W=0.64U L=0.12U M=1 
X8 VDD C Y VDD LPPFET W=1.14U L=0.12U M=1 
X9 VDD B Y VDD LPPFET W=1.14U L=0.12U M=1 
.ENDS NAND3BX2TS 

**** 
*.SUBCKT NAND3BX4TS Y AN B C 
.SUBCKT NAND3BX4TS Y AN B C VSS VDD
X0 VDD AN nmin1 VDD LPPFET W=1.2U L=0.12U M=1 
X1 nmin1 AN VSS VSS LPNFET W=0.86U L=0.12U M=1 
X10 Y nmin1 hnet13 VSS LPNFET W=0.88U L=0.12U M=1 
X11 VDD C Y VDD LPPFET W=2.28U L=0.12U M=1 
X12 VDD B Y VDD LPPFET W=2.28U L=0.12U M=1 
X13 VDD nmin1 Y VDD LPPFET W=2.28U L=0.12U M=1 
X2 hnet20 C VSS VSS LPNFET W=0.88U L=0.12U M=1 
X3 hnet12 B hnet20 VSS LPNFET W=0.88U L=0.12U M=1 
X4 Y nmin1 hnet12 VSS LPNFET W=0.88U L=0.12U M=1 
X5 hnet21 C VSS VSS LPNFET W=0.88U L=0.12U M=1 
X6 hnet16 B hnet21 VSS LPNFET W=0.88U L=0.12U M=1 
X7 Y nmin1 hnet16 VSS LPNFET W=0.88U L=0.12U M=1 
X8 hnet15 C VSS VSS LPNFET W=0.88U L=0.12U M=1 
X9 hnet13 B hnet15 VSS LPNFET W=0.88U L=0.12U M=1 
.ENDS NAND3BX4TS 

**** 
*.SUBCKT NAND3BXLTS Y AN B C 
.SUBCKT NAND3BXLTS Y AN B C VSS VDD
X0 VDD AN nmin1 VDD LPPFET W=0.28U L=0.12U M=1 
X1 nmin1 AN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 hnet17 C VSS VSS LPNFET W=0.48U L=0.12U M=1 
X3 hnet12 B hnet17 VSS LPNFET W=0.48U L=0.12U M=1 
X4 Y nmin1 hnet12 VSS LPNFET W=0.48U L=0.12U M=1 
X5 VDD C Y VDD LPPFET W=0.42U L=0.12U M=1 
X6 VDD B Y VDD LPPFET W=0.42U L=0.12U M=1 
X7 VDD nmin1 Y VDD LPPFET W=0.42U L=0.12U M=1 
.ENDS NAND3BXLTS 

**** 
*.SUBCKT NAND3X1TS Y A B C 
.SUBCKT NAND3X1TS Y A B C VSS VDD
X0 hnet14 C VSS VSS LPNFET W=0.72U L=0.12U M=1 
X1 hnet7 B hnet14 VSS LPNFET W=0.72U L=0.12U M=1 
X2 Y A hnet7 VSS LPNFET W=0.72U L=0.12U M=1 
X3 VDD C Y VDD LPPFET W=0.64U L=0.12U M=1 
X4 VDD B Y VDD LPPFET W=0.64U L=0.12U M=1 
X5 VDD A Y VDD LPPFET W=0.64U L=0.12U M=1 
.ENDS NAND3X1TS 

**** 
*.SUBCKT NAND3X2TS Y A B C 
.SUBCKT NAND3X2TS Y A B C VSS VDD
X0 hnet15 C VSS VSS LPNFET W=0.66U L=0.12U M=1 
X1 hnet7 B hnet15 VSS LPNFET W=0.66U L=0.12U M=1 
X2 Y A hnet7 VSS LPNFET W=0.66U L=0.12U M=1 
X3 hnet16 C VSS VSS LPNFET W=0.66U L=0.12U M=1 
X4 hnet10 B hnet16 VSS LPNFET W=0.66U L=0.12U M=1 
X5 Y A hnet10 VSS LPNFET W=0.66U L=0.12U M=1 
X6 VDD C Y VDD LPPFET W=1.26U L=0.12U M=1 
X7 VDD B Y VDD LPPFET W=1.26U L=0.12U M=1 
X8 VDD A Y VDD LPPFET W=1.26U L=0.12U M=1 
.ENDS NAND3X2TS 

**** 
*.SUBCKT NAND3X4TS Y A B C 
.SUBCKT NAND3X4TS Y A B C VSS VDD
X0 hnet16 C VSS VSS LPNFET W=0.88U L=0.12U M=1 
X1 hnet7 B hnet16 VSS LPNFET W=0.88U L=0.12U M=1 
X10 VDD B Y VDD LPPFET W=2.42U L=0.12U M=1 
X11 VDD A Y VDD LPPFET W=2.42U L=0.12U M=1 
X2 Y A hnet7 VSS LPNFET W=0.88U L=0.12U M=1 
X3 hnet18 C VSS VSS LPNFET W=0.88U L=0.12U M=1 
X4 hnet12 B hnet18 VSS LPNFET W=0.88U L=0.12U M=1 
X5 Y A hnet12 VSS LPNFET W=0.88U L=0.12U M=1 
X6 hnet11 C VSS VSS LPNFET W=0.88U L=0.12U M=1 
X7 hnet8 B hnet11 VSS LPNFET W=0.88U L=0.12U M=1 
X8 Y A hnet8 VSS LPNFET W=0.88U L=0.12U M=1 
X9 VDD C Y VDD LPPFET W=2.42U L=0.12U M=1 
.ENDS NAND3X4TS 

**** 
*.SUBCKT NAND3X6TS Y A B C 
.SUBCKT NAND3X6TS Y A B C VSS VDD
X0 hnet7 C VSS VSS LPNFET W=0.88U L=0.12U M=1 
X1 hnet8 B hnet7 VSS LPNFET W=0.88U L=0.12U M=1 
X10 hnet9 B hnet11 VSS LPNFET W=0.88U L=0.12U M=1 
X11 Y A hnet9 VSS LPNFET W=0.88U L=0.12U M=1 
X12 VDD C Y VDD LPPFET W=3.84U L=0.12U M=1 
X13 VDD B Y VDD LPPFET W=3.84U L=0.12U M=1 
X14 VDD A Y VDD LPPFET W=3.84U L=0.12U M=1 
X2 Y A hnet8 VSS LPNFET W=0.88U L=0.12U M=1 
X3 hnet19 C VSS VSS LPNFET W=0.88U L=0.12U M=1 
X4 hnet20 B hnet19 VSS LPNFET W=0.88U L=0.12U M=1 
X5 Y A hnet20 VSS LPNFET W=0.88U L=0.12U M=1 
X6 hnet14 C VSS VSS LPNFET W=0.88U L=0.12U M=1 
X7 hnet10 B hnet14 VSS LPNFET W=0.88U L=0.12U M=1 
X8 Y A hnet10 VSS LPNFET W=0.88U L=0.12U M=1 
X9 hnet11 C VSS VSS LPNFET W=0.88U L=0.12U M=1 
.ENDS NAND3X6TS 

**** 
*.SUBCKT NAND3X8TS Y A B C 
.SUBCKT NAND3X8TS Y A B C VSS VDD
X0 hnet21 C VSS VSS LPNFET W=0.86U L=0.12U M=1 
X1 hnet8 B hnet21 VSS LPNFET W=0.86U L=0.12U M=1 
X10 hnet7 B hnet10 VSS LPNFET W=0.86U L=0.12U M=1 
X11 Y A hnet7 VSS LPNFET W=0.86U L=0.12U M=1 
X12 hnet23 C VSS VSS LPNFET W=0.86U L=0.12U M=1 
X13 hnet22 B hnet23 VSS LPNFET W=0.86U L=0.12U M=1 
X14 Y A hnet22 VSS LPNFET W=0.86U L=0.12U M=1 
X15 hnet13 C VSS VSS LPNFET W=0.86U L=0.12U M=1 
X16 hnet11 B hnet13 VSS LPNFET W=0.86U L=0.12U M=1 
X17 Y A hnet11 VSS LPNFET W=0.86U L=0.12U M=1 
X18 VDD C Y VDD LPPFET W=4.84U L=0.12U M=1 
X19 VDD B Y VDD LPPFET W=4.84U L=0.12U M=1 
X2 Y A hnet8 VSS LPNFET W=0.86U L=0.12U M=1 
X20 VDD A Y VDD LPPFET W=4.84U L=0.12U M=1 
X3 hnet24 C VSS VSS LPNFET W=0.86U L=0.12U M=1 
X4 hnet16 B hnet24 VSS LPNFET W=0.86U L=0.12U M=1 
X5 Y A hnet16 VSS LPNFET W=0.86U L=0.12U M=1 
X6 hnet15 C VSS VSS LPNFET W=0.86U L=0.12U M=1 
X7 hnet9 B hnet15 VSS LPNFET W=0.86U L=0.12U M=1 
X8 Y A hnet9 VSS LPNFET W=0.86U L=0.12U M=1 
X9 hnet10 C VSS VSS LPNFET W=0.86U L=0.12U M=1 
.ENDS NAND3X8TS 

**** 
*.SUBCKT NAND3XLTS Y A B C 
.SUBCKT NAND3XLTS Y A B C VSS VDD
X0 hnet14 C VSS VSS LPNFET W=0.48U L=0.12U M=1 
X1 hnet7 B hnet14 VSS LPNFET W=0.48U L=0.12U M=1 
X2 Y A hnet7 VSS LPNFET W=0.48U L=0.12U M=1 
X3 VDD C Y VDD LPPFET W=0.42U L=0.12U M=1 
X4 VDD B Y VDD LPPFET W=0.42U L=0.12U M=1 
X5 VDD A Y VDD LPPFET W=0.42U L=0.12U M=1 
.ENDS NAND3XLTS 

**** 
*.SUBCKT NAND4BBX1TS Y AN BN C D 
.SUBCKT NAND4BBX1TS Y AN BN C D VSS VDD
X0 VDD BN nmin2 VDD LPPFET W=0.34U L=0.12U M=1 
X1 nmin2 BN VSS VSS LPNFET W=0.24U L=0.12U M=1 
X10 VDD nmin2 Y VDD LPPFET W=0.64U L=0.12U M=1 
X11 VDD nmin1 Y VDD LPPFET W=0.64U L=0.12U M=1 
X2 VDD AN nmin1 VDD LPPFET W=0.34U L=0.12U M=1 
X3 nmin1 AN VSS VSS LPNFET W=0.24U L=0.12U M=1 
X4 hnet19 D VSS VSS LPNFET W=0.78U L=0.12U M=1 
X5 hnet18 C hnet19 VSS LPNFET W=0.78U L=0.12U M=1 
X6 hnet20 nmin2 hnet18 VSS LPNFET W=0.78U L=0.12U M=1 
X7 Y nmin1 hnet20 VSS LPNFET W=0.78U L=0.12U M=1 
X8 VDD D Y VDD LPPFET W=0.64U L=0.12U M=1 
X9 VDD C Y VDD LPPFET W=0.64U L=0.12U M=1 
.ENDS NAND4BBX1TS 

**** 
*.SUBCKT NAND4BBX2TS Y AN BN C D 
.SUBCKT NAND4BBX2TS Y AN BN C D VSS VDD
X0 VDD BN nmin2 VDD LPPFET W=0.66U L=0.12U M=1 
X1 nmin2 BN VSS VSS LPNFET W=0.48U L=0.12U M=1 
X10 hnet22 nmin2 hnet27 VSS LPNFET W=0.8U L=0.12U M=1 
X11 Y nmin1 hnet22 VSS LPNFET W=0.8U L=0.12U M=1 
X12 VDD D Y VDD LPPFET W=1.24U L=0.12U M=1 
X13 VDD C Y VDD LPPFET W=1.24U L=0.12U M=1 
X14 VDD nmin2 Y VDD LPPFET W=1.24U L=0.12U M=1 
X15 VDD nmin1 Y VDD LPPFET W=1.24U L=0.12U M=1 
X2 VDD AN nmin1 VDD LPPFET W=0.66U L=0.12U M=1 
X3 nmin1 AN VSS VSS LPNFET W=0.48U L=0.12U M=1 
X4 hnet18 D VSS VSS LPNFET W=0.8U L=0.12U M=1 
X5 hnet19 C hnet18 VSS LPNFET W=0.8U L=0.12U M=1 
X6 hnet20 nmin2 hnet19 VSS LPNFET W=0.8U L=0.12U M=1 
X7 Y nmin1 hnet20 VSS LPNFET W=0.8U L=0.12U M=1 
X8 hnet23 D VSS VSS LPNFET W=0.8U L=0.12U M=1 
X9 hnet27 C hnet23 VSS LPNFET W=0.8U L=0.12U M=1 
.ENDS NAND4BBX2TS 

**** 
*.SUBCKT NAND4BBX4TS Y AN BN C D 
.SUBCKT NAND4BBX4TS Y AN BN C D VSS VDD
X0 VDD BN nmin2 VDD LPPFET W=1.3U L=0.12U M=1 
X1 nmin2 BN VSS VSS LPNFET W=0.92U L=0.12U M=1 
X10 hnet26 nmin2 hnet30 VSS LPNFET W=0.76U L=0.12U M=1 
X11 Y nmin1 hnet26 VSS LPNFET W=0.76U L=0.12U M=1 
X12 hnet24 D VSS VSS LPNFET W=0.76U L=0.12U M=1 
X13 hnet21 C hnet24 VSS LPNFET W=0.76U L=0.12U M=1 
X14 hnet18 nmin2 hnet21 VSS LPNFET W=0.76U L=0.12U M=1 
X15 Y nmin1 hnet18 VSS LPNFET W=0.76U L=0.12U M=1 
X16 hnet33 D VSS VSS LPNFET W=0.76U L=0.12U M=1 
X17 hnet27 C hnet33 VSS LPNFET W=0.76U L=0.12U M=1 
X18 hnet23 nmin2 hnet27 VSS LPNFET W=0.76U L=0.12U M=1 
X19 Y nmin1 hnet23 VSS LPNFET W=0.76U L=0.12U M=1 
X2 VDD AN nmin1 VDD LPPFET W=1.3U L=0.12U M=1 
X20 VDD D Y VDD LPPFET W=2.54U L=0.12U M=1 
X21 VDD C Y VDD LPPFET W=2.54U L=0.12U M=1 
X22 VDD nmin2 Y VDD LPPFET W=2.54U L=0.12U M=1 
X23 VDD nmin1 Y VDD LPPFET W=2.54U L=0.12U M=1 
X3 nmin1 AN VSS VSS LPNFET W=0.92U L=0.12U M=1 
X4 hnet20 D VSS VSS LPNFET W=0.76U L=0.12U M=1 
X5 hnet19 C hnet20 VSS LPNFET W=0.76U L=0.12U M=1 
X6 hnet22 nmin2 hnet19 VSS LPNFET W=0.76U L=0.12U M=1 
X7 Y nmin1 hnet22 VSS LPNFET W=0.76U L=0.12U M=1 
X8 hnet28 D VSS VSS LPNFET W=0.76U L=0.12U M=1 
X9 hnet30 C hnet28 VSS LPNFET W=0.76U L=0.12U M=1 
.ENDS NAND4BBX4TS 

**** 
*.SUBCKT NAND4BBXLTS Y AN BN C D 
.SUBCKT NAND4BBXLTS Y AN BN C D VSS VDD
X0 VDD BN nmin2 VDD LPPFET W=0.28U L=0.12U M=1 
X1 nmin2 BN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X10 VDD nmin2 Y VDD LPPFET W=0.42U L=0.12U M=1 
X11 VDD nmin1 Y VDD LPPFET W=0.42U L=0.12U M=1 
X2 VDD AN nmin1 VDD LPPFET W=0.28U L=0.12U M=1 
X3 nmin1 AN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X4 hnet19 D VSS VSS LPNFET W=0.52U L=0.12U M=1 
X5 hnet18 C hnet19 VSS LPNFET W=0.52U L=0.12U M=1 
X6 hnet20 nmin2 hnet18 VSS LPNFET W=0.52U L=0.12U M=1 
X7 Y nmin1 hnet20 VSS LPNFET W=0.52U L=0.12U M=1 
X8 VDD D Y VDD LPPFET W=0.42U L=0.12U M=1 
X9 VDD C Y VDD LPPFET W=0.42U L=0.12U M=1 
.ENDS NAND4BBXLTS 

**** 
*.SUBCKT NAND4BX1TS Y AN B C D 
.SUBCKT NAND4BX1TS Y AN B C D VSS VDD
X0 VDD AN nmin1 VDD LPPFET W=0.34U L=0.12U M=1 
X1 nmin1 AN VSS VSS LPNFET W=0.24U L=0.12U M=1 
X2 hnet14 D VSS VSS LPNFET W=0.78U L=0.12U M=1 
X3 hnet13 C hnet14 VSS LPNFET W=0.78U L=0.12U M=1 
X4 hnet15 B hnet13 VSS LPNFET W=0.78U L=0.12U M=1 
X5 Y nmin1 hnet15 VSS LPNFET W=0.78U L=0.12U M=1 
X6 VDD D Y VDD LPPFET W=0.64U L=0.12U M=1 
X7 VDD C Y VDD LPPFET W=0.64U L=0.12U M=1 
X8 VDD B Y VDD LPPFET W=0.64U L=0.12U M=1 
X9 VDD nmin1 Y VDD LPPFET W=0.64U L=0.12U M=1 
.ENDS NAND4BX1TS 

**** 
*.SUBCKT NAND4BX2TS Y AN B C D 
.SUBCKT NAND4BX2TS Y AN B C D VSS VDD
X0 VDD AN nmin1 VDD LPPFET W=0.66U L=0.12U M=1 
X1 nmin1 AN VSS VSS LPNFET W=0.48U L=0.12U M=1 
X10 VDD D Y VDD LPPFET W=1.22U L=0.12U M=1 
X11 VDD C Y VDD LPPFET W=1.22U L=0.12U M=1 
X12 VDD B Y VDD LPPFET W=1.22U L=0.12U M=1 
X13 VDD nmin1 Y VDD LPPFET W=1.22U L=0.12U M=1 
X2 hnet13 D VSS VSS LPNFET W=0.8U L=0.12U M=1 
X3 hnet14 C hnet13 VSS LPNFET W=0.8U L=0.12U M=1 
X4 hnet15 B hnet14 VSS LPNFET W=0.8U L=0.12U M=1 
X5 Y nmin1 hnet15 VSS LPNFET W=0.8U L=0.12U M=1 
X6 hnet18 D VSS VSS LPNFET W=0.8U L=0.12U M=1 
X7 hnet22 C hnet18 VSS LPNFET W=0.8U L=0.12U M=1 
X8 hnet17 B hnet22 VSS LPNFET W=0.8U L=0.12U M=1 
X9 Y nmin1 hnet17 VSS LPNFET W=0.8U L=0.12U M=1 
.ENDS NAND4BX2TS 

**** 
*.SUBCKT NAND4BX4TS Y AN B C D 
.SUBCKT NAND4BX4TS Y AN B C D VSS VDD
X0 VDD AN nmin1 VDD LPPFET W=1.3U L=0.12U M=1 
X1 nmin1 AN VSS VSS LPNFET W=0.92U L=0.12U M=1 
X10 hnet19 D VSS VSS LPNFET W=0.74U L=0.12U M=1 
X11 hnet16 C hnet19 VSS LPNFET W=0.74U L=0.12U M=1 
X12 hnet13 B hnet16 VSS LPNFET W=0.74U L=0.12U M=1 
X13 Y nmin1 hnet13 VSS LPNFET W=0.74U L=0.12U M=1 
X14 hnet28 D VSS VSS LPNFET W=0.74U L=0.12U M=1 
X15 hnet22 C hnet28 VSS LPNFET W=0.74U L=0.12U M=1 
X16 hnet18 B hnet22 VSS LPNFET W=0.74U L=0.12U M=1 
X17 Y nmin1 hnet18 VSS LPNFET W=0.74U L=0.12U M=1 
X18 VDD D Y VDD LPPFET W=2.54U L=0.12U M=1 
X19 VDD C Y VDD LPPFET W=2.54U L=0.12U M=1 
X2 hnet15 D VSS VSS LPNFET W=0.74U L=0.12U M=1 
X20 VDD B Y VDD LPPFET W=2.54U L=0.12U M=1 
X21 VDD nmin1 Y VDD LPPFET W=2.54U L=0.12U M=1 
X3 hnet14 C hnet15 VSS LPNFET W=0.74U L=0.12U M=1 
X4 hnet17 B hnet14 VSS LPNFET W=0.74U L=0.12U M=1 
X5 Y nmin1 hnet17 VSS LPNFET W=0.74U L=0.12U M=1 
X6 hnet23 D VSS VSS LPNFET W=0.74U L=0.12U M=1 
X7 hnet25 C hnet23 VSS LPNFET W=0.74U L=0.12U M=1 
X8 hnet21 B hnet25 VSS LPNFET W=0.74U L=0.12U M=1 
X9 Y nmin1 hnet21 VSS LPNFET W=0.74U L=0.12U M=1 
.ENDS NAND4BX4TS 

**** 
*.SUBCKT NAND4BXLTS Y AN B C D 
.SUBCKT NAND4BXLTS Y AN B C D VSS VDD
X0 VDD AN nmin1 VDD LPPFET W=0.28U L=0.12U M=1 
X1 nmin1 AN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 hnet14 D VSS VSS LPNFET W=0.52U L=0.12U M=1 
X3 hnet13 C hnet14 VSS LPNFET W=0.52U L=0.12U M=1 
X4 hnet15 B hnet13 VSS LPNFET W=0.52U L=0.12U M=1 
X5 Y nmin1 hnet15 VSS LPNFET W=0.52U L=0.12U M=1 
X6 VDD D Y VDD LPPFET W=0.42U L=0.12U M=1 
X7 VDD C Y VDD LPPFET W=0.42U L=0.12U M=1 
X8 VDD B Y VDD LPPFET W=0.42U L=0.12U M=1 
X9 VDD nmin1 Y VDD LPPFET W=0.42U L=0.12U M=1 
.ENDS NAND4BXLTS 

**** 
*.SUBCKT NAND4X1TS Y A B C D 
.SUBCKT NAND4X1TS Y A B C D VSS VDD
X0 hnet9 D VSS VSS LPNFET W=0.78U L=0.12U M=1 
X1 hnet8 C hnet9 VSS LPNFET W=0.78U L=0.12U M=1 
X2 hnet10 B hnet8 VSS LPNFET W=0.78U L=0.12U M=1 
X3 Y A hnet10 VSS LPNFET W=0.78U L=0.12U M=1 
X4 VDD D Y VDD LPPFET W=0.64U L=0.12U M=1 
X5 VDD C Y VDD LPPFET W=0.64U L=0.12U M=1 
X6 VDD B Y VDD LPPFET W=0.64U L=0.12U M=1 
X7 VDD A Y VDD LPPFET W=0.64U L=0.12U M=1 
.ENDS NAND4X1TS 

**** 
*.SUBCKT NAND4X2TS Y A B C D 
.SUBCKT NAND4X2TS Y A B C D VSS VDD
X0 hnet8 D VSS VSS LPNFET W=0.78U L=0.12U M=1 
X1 hnet9 C hnet8 VSS LPNFET W=0.78U L=0.12U M=1 
X10 VDD B Y VDD LPPFET W=1.18U L=0.12U M=1 
X11 VDD A Y VDD LPPFET W=1.18U L=0.12U M=1 
X2 hnet10 B hnet9 VSS LPNFET W=0.78U L=0.12U M=1 
X3 Y A hnet10 VSS LPNFET W=0.78U L=0.12U M=1 
X4 hnet14 D VSS VSS LPNFET W=0.78U L=0.12U M=1 
X5 hnet19 C hnet14 VSS LPNFET W=0.78U L=0.12U M=1 
X6 hnet12 B hnet19 VSS LPNFET W=0.78U L=0.12U M=1 
X7 Y A hnet12 VSS LPNFET W=0.78U L=0.12U M=1 
X8 VDD D Y VDD LPPFET W=1.18U L=0.12U M=1 
X9 VDD C Y VDD LPPFET W=1.18U L=0.12U M=1 
.ENDS NAND4X2TS 

**** 
*.SUBCKT NAND4X4TS Y A B C D 
.SUBCKT NAND4X4TS Y A B C D VSS VDD
X0 hnet10 D VSS VSS LPNFET W=0.78U L=0.12U M=1 
X1 hnet9 C hnet10 VSS LPNFET W=0.78U L=0.12U M=1 
X10 hnet8 B hnet11 VSS LPNFET W=0.78U L=0.12U M=1 
X11 Y A hnet8 VSS LPNFET W=0.78U L=0.12U M=1 
X12 hnet25 D VSS VSS LPNFET W=0.78U L=0.12U M=1 
X13 hnet17 C hnet25 VSS LPNFET W=0.78U L=0.12U M=1 
X14 hnet13 B hnet17 VSS LPNFET W=0.78U L=0.12U M=1 
X15 Y A hnet13 VSS LPNFET W=0.78U L=0.12U M=1 
X16 VDD D Y VDD LPPFET W=2.44U L=0.12U M=1 
X17 VDD C Y VDD LPPFET W=2.44U L=0.12U M=1 
X18 VDD B Y VDD LPPFET W=2.44U L=0.12U M=1 
X19 VDD A Y VDD LPPFET W=2.44U L=0.12U M=1 
X2 hnet12 B hnet9 VSS LPNFET W=0.78U L=0.12U M=1 
X3 Y A hnet12 VSS LPNFET W=0.78U L=0.12U M=1 
X4 hnet19 D VSS VSS LPNFET W=0.78U L=0.12U M=1 
X5 hnet21 C hnet19 VSS LPNFET W=0.78U L=0.12U M=1 
X6 hnet16 B hnet21 VSS LPNFET W=0.78U L=0.12U M=1 
X7 Y A hnet16 VSS LPNFET W=0.78U L=0.12U M=1 
X8 hnet14 D VSS VSS LPNFET W=0.78U L=0.12U M=1 
X9 hnet11 C hnet14 VSS LPNFET W=0.78U L=0.12U M=1 
.ENDS NAND4X4TS 

**** 
*.SUBCKT NAND4X6TS Y A B C D 
.SUBCKT NAND4X6TS Y A B C D VSS VDD
X0 hnet28 D VSS VSS LPNFET W=0.82U L=0.12U M=1 
X1 hnet8 C hnet28 VSS LPNFET W=0.82U L=0.12U M=1 
X10 hnet24 B hnet12 VSS LPNFET W=0.82U L=0.12U M=1 
X11 Y A hnet24 VSS LPNFET W=0.82U L=0.12U M=1 
X12 hnet25 D VSS VSS LPNFET W=0.82U L=0.12U M=1 
X13 hnet16 C hnet25 VSS LPNFET W=0.82U L=0.12U M=1 
X14 hnet13 B hnet16 VSS LPNFET W=0.82U L=0.12U M=1 
X15 Y A hnet13 VSS LPNFET W=0.82U L=0.12U M=1 
X16 hnet9 D VSS VSS LPNFET W=0.82U L=0.12U M=1 
X17 hnet29 C hnet9 VSS LPNFET W=0.82U L=0.12U M=1 
X18 hnet26 B hnet29 VSS LPNFET W=0.82U L=0.12U M=1 
X19 Y A hnet26 VSS LPNFET W=0.82U L=0.12U M=1 
X2 hnet11 B hnet8 VSS LPNFET W=0.82U L=0.12U M=1 
X20 VDD D Y VDD LPPFET W=3.68U L=0.12U M=1 
X21 VDD C Y VDD LPPFET W=3.68U L=0.12U M=1 
X22 VDD B Y VDD LPPFET W=3.68U L=0.12U M=1 
X23 VDD A Y VDD LPPFET W=3.68U L=0.12U M=1 
X3 Y A hnet11 VSS LPNFET W=0.82U L=0.12U M=1 
X4 hnet18 D VSS VSS LPNFET W=0.82U L=0.12U M=1 
X5 hnet20 C hnet18 VSS LPNFET W=0.82U L=0.12U M=1 
X6 hnet15 B hnet20 VSS LPNFET W=0.82U L=0.12U M=1 
X7 Y A hnet15 VSS LPNFET W=0.82U L=0.12U M=1 
X8 hnet10 D VSS VSS LPNFET W=0.82U L=0.12U M=1 
X9 hnet12 C hnet10 VSS LPNFET W=0.82U L=0.12U M=1 
.ENDS NAND4X6TS 

**** 
*.SUBCKT NAND4X8TS Y A B C D 
.SUBCKT NAND4X8TS Y A B C D VSS VDD
X0 hnet11 D VSS VSS LPNFET W=0.86U L=0.12U M=1 
X1 hnet13 C hnet11 VSS LPNFET W=0.86U L=0.12U M=1 
X10 hnet26 B hnet25 VSS LPNFET W=0.86U L=0.12U M=1 
X11 Y A hnet26 VSS LPNFET W=0.86U L=0.12U M=1 
X12 hnet15 D VSS VSS LPNFET W=0.86U L=0.12U M=1 
X13 hnet14 C hnet15 VSS LPNFET W=0.86U L=0.12U M=1 
X14 hnet31 B hnet14 VSS LPNFET W=0.86U L=0.12U M=1 
X15 Y A hnet31 VSS LPNFET W=0.86U L=0.12U M=1 
X16 hnet30 D VSS VSS LPNFET W=0.86U L=0.12U M=1 
X17 hnet20 C hnet30 VSS LPNFET W=0.86U L=0.12U M=1 
X18 hnet12 B hnet20 VSS LPNFET W=0.86U L=0.12U M=1 
X19 Y A hnet12 VSS LPNFET W=0.86U L=0.12U M=1 
X2 hnet23 B hnet13 VSS LPNFET W=0.86U L=0.12U M=1 
X20 hnet9 D VSS VSS LPNFET W=0.86U L=0.12U M=1 
X21 hnet35 C hnet9 VSS LPNFET W=0.86U L=0.12U M=1 
X22 hnet32 B hnet35 VSS LPNFET W=0.86U L=0.12U M=1 
X23 Y A hnet32 VSS LPNFET W=0.86U L=0.12U M=1 
X24 hnet17 D VSS VSS LPNFET W=0.86U L=0.12U M=1 
X25 hnet16 C hnet17 VSS LPNFET W=0.86U L=0.12U M=1 
X26 hnet19 B hnet16 VSS LPNFET W=0.86U L=0.12U M=1 
X27 Y A hnet19 VSS LPNFET W=0.86U L=0.12U M=1 
X28 VDD D Y VDD LPPFET W=4.72U L=0.12U M=1 
X29 VDD C Y VDD LPPFET W=4.72U L=0.12U M=1 
X3 Y A hnet23 VSS LPNFET W=0.86U L=0.12U M=1 
X30 VDD B Y VDD LPPFET W=4.72U L=0.12U M=1 
X31 VDD A Y VDD LPPFET W=4.72U L=0.12U M=1 
X4 hnet34 D VSS VSS LPNFET W=0.86U L=0.12U M=1 
X5 hnet8 C hnet34 VSS LPNFET W=0.86U L=0.12U M=1 
X6 hnet10 B hnet8 VSS LPNFET W=0.86U L=0.12U M=1 
X7 Y A hnet10 VSS LPNFET W=0.86U L=0.12U M=1 
X8 hnet22 D VSS VSS LPNFET W=0.86U L=0.12U M=1 
X9 hnet25 C hnet22 VSS LPNFET W=0.86U L=0.12U M=1 
.ENDS NAND4X8TS 

**** 
*.SUBCKT NAND4XLTS Y A B C D 
.SUBCKT NAND4XLTS Y A B C D VSS VDD
X0 hnet9 D VSS VSS LPNFET W=0.52U L=0.12U M=1 
X1 hnet8 C hnet9 VSS LPNFET W=0.52U L=0.12U M=1 
X2 hnet10 B hnet8 VSS LPNFET W=0.52U L=0.12U M=1 
X3 Y A hnet10 VSS LPNFET W=0.52U L=0.12U M=1 
X4 VDD D Y VDD LPPFET W=0.42U L=0.12U M=1 
X5 VDD C Y VDD LPPFET W=0.42U L=0.12U M=1 
X6 VDD B Y VDD LPPFET W=0.42U L=0.12U M=1 
X7 VDD A Y VDD LPPFET W=0.42U L=0.12U M=1 
.ENDS NAND4XLTS 

**** 
*.SUBCKT NOR2BX1TS Y AN B 
.SUBCKT NOR2BX1TS Y AN B VSS VDD
X0 VDD AN nmin1 VDD LPPFET W=0.3U L=0.12U M=1 
X1 nmin1 AN VSS VSS LPNFET W=0.22U L=0.12U M=1 
X2 Y B VSS VSS LPNFET W=0.46U L=0.12U M=1 
X3 Y nmin1 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X4 VDD B hnet12 VDD LPPFET W=0.84U L=0.12U M=1 
X5 hnet12 nmin1 Y VDD LPPFET W=0.84U L=0.12U M=1 
.ENDS NOR2BX1TS 

**** 
*.SUBCKT NOR2BX2TS Y AN B 
.SUBCKT NOR2BX2TS Y AN B VSS VDD
X0 VDD AN nmin1 VDD LPPFET W=0.62U L=0.12U M=1 
X1 nmin1 AN VSS VSS LPNFET W=0.44U L=0.12U M=1 
X2 Y B VSS VSS LPNFET W=0.92U L=0.12U M=1 
X3 Y nmin1 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X4 VDD B hnet13 VDD LPPFET W=0.84U L=0.12U M=1 
X5 hnet13 nmin1 Y VDD LPPFET W=0.84U L=0.12U M=1 
X6 VDD B hnet11 VDD LPPFET W=0.84U L=0.12U M=1 
X7 hnet11 nmin1 Y VDD LPPFET W=0.84U L=0.12U M=1 
.ENDS NOR2BX2TS 

**** 
*.SUBCKT NOR2BX4TS Y AN B 
.SUBCKT NOR2BX4TS Y AN B VSS VDD
X0 VDD AN nmin1 VDD LPPFET W=1.2U L=0.12U M=1 
X1 nmin1 AN VSS VSS LPNFET W=0.86U L=0.12U M=1 
X2 Y B VSS VSS LPNFET W=1.84U L=0.12U M=1 
X3 Y nmin1 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X4 VDD B hnet13 VDD LPPFET W=1.04U L=0.12U M=1 
X5 hnet13 nmin1 Y VDD LPPFET W=1.04U L=0.12U M=1 
X6 VDD B hnet11 VDD LPPFET W=1.04U L=0.12U M=1 
X7 hnet11 nmin1 Y VDD LPPFET W=1.04U L=0.12U M=1 
X8 VDD B hnet14 VDD LPPFET W=1.04U L=0.12U M=1 
X9 hnet14 nmin1 Y VDD LPPFET W=1.04U L=0.12U M=1 
.ENDS NOR2BX4TS 

**** 
*.SUBCKT NOR2BXLTS Y AN B 
.SUBCKT NOR2BXLTS Y AN B VSS VDD
X0 VDD AN nmin1 VDD LPPFET W=0.28U L=0.12U M=1 
X1 nmin1 AN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 Y B VSS VSS LPNFET W=0.24U L=0.12U M=1 
X3 Y nmin1 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X4 VDD B hnet12 VDD LPPFET W=0.44U L=0.12U M=1 
X5 hnet12 nmin1 Y VDD LPPFET W=0.44U L=0.12U M=1 
.ENDS NOR2BXLTS 

**** 
*.SUBCKT NOR2X1TS Y A B 
.SUBCKT NOR2X1TS Y A B VSS VDD
X0 Y B VSS VSS LPNFET W=0.46U L=0.12U M=1 
X1 Y A VSS VSS LPNFET W=0.46U L=0.12U M=1 
X2 VDD B hnet7 VDD LPPFET W=0.84U L=0.12U M=1 
X3 hnet7 A Y VDD LPPFET W=0.84U L=0.12U M=1 
.ENDS NOR2X1TS 

**** 
*.SUBCKT NOR2X2TS Y A B 
.SUBCKT NOR2X2TS Y A B VSS VDD
X0 Y B VSS VSS LPNFET W=0.92U L=0.12U M=1 
X1 Y A VSS VSS LPNFET W=0.92U L=0.12U M=1 
X2 VDD B hnet8 VDD LPPFET W=0.84U L=0.12U M=1 
X3 hnet8 A Y VDD LPPFET W=0.84U L=0.12U M=1 
X4 VDD B hnet6 VDD LPPFET W=0.84U L=0.12U M=1 
X5 hnet6 A Y VDD LPPFET W=0.84U L=0.12U M=1 
.ENDS NOR2X2TS 

**** 
*.SUBCKT NOR2X4TS Y A B 
.SUBCKT NOR2X4TS Y A B VSS VDD
X0 VDD B net15 VDD LPPFET W=1.12U L=0.12U M=1 
X1 net15 A Y VDD LPPFET W=1.12U L=0.12U M=1 
X2 VDD B net17 VDD LPPFET W=1.12U L=0.12U M=1 
X3 net17 A Y VDD LPPFET W=1.12U L=0.12U M=1 
X4 VDD B net27 VDD LPPFET W=1.06U L=0.12U M=1 
X5 net27 A Y VDD LPPFET W=1.06U L=0.12U M=1 
X6 Y B VSS VSS LPNFET W=1.84U L=0.12U M=1 
X7 Y A VSS VSS LPNFET W=1.84U L=0.12U M=1 
.ENDS NOR2X4TS 

**** 
*.SUBCKT NOR2X6TS Y A B 
.SUBCKT NOR2X6TS Y A B VSS VDD
X0 Y B VSS VSS LPNFET W=2.76U L=0.12U M=1 
X1 Y A VSS VSS LPNFET W=2.76U L=0.12U M=1 
X2 VDD B hnet9 VDD LPPFET W=1.16U L=0.12U M=1 
X3 hnet9 A Y VDD LPPFET W=1.16U L=0.12U M=1 
X4 VDD B hnet6 VDD LPPFET W=1.16U L=0.12U M=1 
X5 hnet6 A Y VDD LPPFET W=1.16U L=0.12U M=1 
X6 VDD B hnet11 VDD LPPFET W=1.16U L=0.12U M=1 
X7 hnet11 A Y VDD LPPFET W=1.16U L=0.12U M=1 
X8 VDD B hnet8 VDD LPPFET W=1.16U L=0.12U M=1 
X9 hnet8 A Y VDD LPPFET W=1.16U L=0.12U M=1 
.ENDS NOR2X6TS 

**** 
*.SUBCKT NOR2X8TS Y A B 
.SUBCKT NOR2X8TS Y A B VSS VDD
X0 Y B VSS VSS LPNFET W=3.44U L=0.12U M=1 
X1 Y A VSS VSS LPNFET W=3.44U L=0.12U M=1 
X10 VDD B hnet6 VDD LPPFET W=1.3U L=0.12U M=1 
X11 hnet6 A Y VDD LPPFET W=1.3U L=0.12U M=1 
X2 VDD B hnet9 VDD LPPFET W=1.3U L=0.12U M=1 
X3 hnet9 A Y VDD LPPFET W=1.3U L=0.12U M=1 
X4 VDD B hnet8 VDD LPPFET W=1.3U L=0.12U M=1 
X5 hnet8 A Y VDD LPPFET W=1.3U L=0.12U M=1 
X6 VDD B hnet12 VDD LPPFET W=1.3U L=0.12U M=1 
X7 hnet12 A Y VDD LPPFET W=1.3U L=0.12U M=1 
X8 VDD B hnet7 VDD LPPFET W=1.3U L=0.12U M=1 
X9 hnet7 A Y VDD LPPFET W=1.3U L=0.12U M=1 
.ENDS NOR2X8TS 

**** 
*.SUBCKT NOR2XLTS Y A B 
.SUBCKT NOR2XLTS Y A B VSS VDD
X0 Y B VSS VSS LPNFET W=0.24U L=0.12U M=1 
X1 Y A VSS VSS LPNFET W=0.24U L=0.12U M=1 
X2 VDD B hnet7 VDD LPPFET W=0.44U L=0.12U M=1 
X3 hnet7 A Y VDD LPPFET W=0.44U L=0.12U M=1 
.ENDS NOR2XLTS 

**** 
*.SUBCKT NOR3BX1TS Y AN B C 
.SUBCKT NOR3BX1TS Y AN B C VSS VDD
X0 VDD AN nmin1 VDD LPPFET W=0.34U L=0.12U M=1 
X1 nmin1 AN VSS VSS LPNFET W=0.24U L=0.12U M=1 
X2 Y C VSS VSS LPNFET W=0.46U L=0.12U M=1 
X3 Y B VSS VSS LPNFET W=0.46U L=0.12U M=1 
X4 Y nmin1 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X5 VDD C hnet17 VDD LPPFET W=1.02U L=0.12U M=1 
X6 hnet17 B hnet16 VDD LPPFET W=1.02U L=0.12U M=1 
X7 hnet16 nmin1 Y VDD LPPFET W=1.02U L=0.12U M=1 
.ENDS NOR3BX1TS 

**** 
*.SUBCKT NOR3BX2TS Y AN B C 
.SUBCKT NOR3BX2TS Y AN B C VSS VDD
X0 VDD AN nmin1 VDD LPPFET W=0.64U L=0.12U M=1 
X1 nmin1 AN VSS VSS LPNFET W=0.5U L=0.12U M=1 
X10 hnet12 nmin1 Y VDD LPPFET W=1.04U L=0.12U M=1 
X2 Y C VSS VSS LPNFET W=0.92U L=0.12U M=1 
X3 Y B VSS VSS LPNFET W=0.92U L=0.12U M=1 
X4 Y nmin1 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X5 VDD C hnet19 VDD LPPFET W=1.04U L=0.12U M=1 
X6 hnet19 B hnet15 VDD LPPFET W=1.04U L=0.12U M=1 
X7 hnet15 nmin1 Y VDD LPPFET W=1.04U L=0.12U M=1 
X8 VDD C hnet14 VDD LPPFET W=1.04U L=0.12U M=1 
X9 hnet14 B hnet12 VDD LPPFET W=1.04U L=0.12U M=1 
.ENDS NOR3BX2TS 

**** 
*.SUBCKT NOR3BX4TS Y AN B C 
.SUBCKT NOR3BX4TS Y AN B C VSS VDD
X0 Y C VSS VSS LPNFET W=1.84U L=0.12U M=1 
X1 Y B VSS VSS LPNFET W=1.84U L=0.12U M=1 
X10 hnet9 B hnet10 VDD LPPFET W=0.88U L=0.12U M=1 
X11 hnet10 nmin1 Y VDD LPPFET W=0.88U L=0.12U M=1 
X12 VDD C hnet18 VDD LPPFET W=0.88U L=0.12U M=1 
X13 hnet18 B hnet21 VDD LPPFET W=0.88U L=0.12U M=1 
X14 hnet21 nmin1 Y VDD LPPFET W=0.88U L=0.12U M=1 
X15 VDD AN nmin1 VDD LPPFET W=1.3U L=0.12U M=1 
X16 nmin1 AN VSS VSS LPNFET W=0.92U L=0.12U M=1 
X2 Y nmin1 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X3 VDD C hnet20 VDD LPPFET W=0.88U L=0.12U M=1 
X4 hnet20 B hnet19 VDD LPPFET W=0.88U L=0.12U M=1 
X5 hnet19 nmin1 Y VDD LPPFET W=0.88U L=0.12U M=1 
X6 VDD C hnet12 VDD LPPFET W=0.88U L=0.12U M=1 
X7 hnet12 B hnet8 VDD LPPFET W=0.88U L=0.12U M=1 
X8 hnet8 nmin1 Y VDD LPPFET W=0.88U L=0.12U M=1 
X9 VDD C hnet9 VDD LPPFET W=0.88U L=0.12U M=1 
.ENDS NOR3BX4TS 

**** 
*.SUBCKT NOR3BXLTS Y AN B C 
.SUBCKT NOR3BXLTS Y AN B C VSS VDD
X0 VDD AN nmin1 VDD LPPFET W=0.28U L=0.12U M=1 
X1 nmin1 AN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 Y C VSS VSS LPNFET W=0.24U L=0.12U M=1 
X3 Y B VSS VSS LPNFET W=0.24U L=0.12U M=1 
X4 Y nmin1 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X5 VDD C hnet17 VDD LPPFET W=0.54U L=0.12U M=1 
X6 hnet17 B hnet16 VDD LPPFET W=0.54U L=0.12U M=1 
X7 hnet16 nmin1 Y VDD LPPFET W=0.54U L=0.12U M=1 
.ENDS NOR3BXLTS 

**** 
*.SUBCKT NOR3X1TS Y A B C 
.SUBCKT NOR3X1TS Y A B C VSS VDD
X0 Y C VSS VSS LPNFET W=0.46U L=0.12U M=1 
X1 Y B VSS VSS LPNFET W=0.46U L=0.12U M=1 
X2 Y A VSS VSS LPNFET W=0.46U L=0.12U M=1 
X3 VDD C hnet14 VDD LPPFET W=1.02U L=0.12U M=1 
X4 hnet14 B hnet13 VDD LPPFET W=1.02U L=0.12U M=1 
X5 hnet13 A Y VDD LPPFET W=1.02U L=0.12U M=1 
.ENDS NOR3X1TS 

**** 
*.SUBCKT NOR3X2TS Y A B C 
.SUBCKT NOR3X2TS Y A B C VSS VDD
X0 Y C VSS VSS LPNFET W=0.84U L=0.12U M=1 
X1 Y B VSS VSS LPNFET W=0.84U L=0.12U M=1 
X2 Y A VSS VSS LPNFET W=0.84U L=0.12U M=1 
X3 VDD C hnet16 VDD LPPFET W=0.94U L=0.12U M=1 
X4 hnet16 B hnet11 VDD LPPFET W=0.94U L=0.12U M=1 
X5 hnet11 A Y VDD LPPFET W=0.94U L=0.12U M=1 
X6 VDD C hnet9 VDD LPPFET W=0.94U L=0.12U M=1 
X7 hnet9 B hnet7 VDD LPPFET W=0.94U L=0.12U M=1 
X8 hnet7 A Y VDD LPPFET W=0.94U L=0.12U M=1 
.ENDS NOR3X2TS 

**** 
*.SUBCKT NOR3X4TS Y A B C 
.SUBCKT NOR3X4TS Y A B C VSS VDD
X0 Y C VSS VSS LPNFET W=1.84U L=0.12U M=1 
X1 Y B VSS VSS LPNFET W=1.84U L=0.12U M=1 
X10 hnet8 B hnet9 VDD LPPFET W=0.98U L=0.12U M=1 
X11 hnet9 A Y VDD LPPFET W=0.98U L=0.12U M=1 
X12 VDD C hnet17 VDD LPPFET W=0.98U L=0.12U M=1 
X13 hnet17 B hnet20 VDD LPPFET W=0.98U L=0.12U M=1 
X14 hnet20 A Y VDD LPPFET W=0.98U L=0.12U M=1 
X2 Y A VSS VSS LPNFET W=1.84U L=0.12U M=1 
X3 VDD C hnet19 VDD LPPFET W=0.98U L=0.12U M=1 
X4 hnet19 B hnet18 VDD LPPFET W=0.98U L=0.12U M=1 
X5 hnet18 A Y VDD LPPFET W=0.98U L=0.12U M=1 
X6 VDD C hnet11 VDD LPPFET W=0.98U L=0.12U M=1 
X7 hnet11 B hnet7 VDD LPPFET W=0.98U L=0.12U M=1 
X8 hnet7 A Y VDD LPPFET W=0.98U L=0.12U M=1 
X9 VDD C hnet8 VDD LPPFET W=0.98U L=0.12U M=1 
.ENDS NOR3X4TS 

**** 
*.SUBCKT NOR3X6TS Y A B C 
.SUBCKT NOR3X6TS Y A B C VSS VDD
X0 Y C VSS VSS LPNFET W=2.76U L=0.12U M=1 
X1 Y B VSS VSS LPNFET W=2.76U L=0.12U M=1 
X10 hnet7 B hnet18 VDD LPPFET W=1.24U L=0.12U M=1 
X11 hnet18 A Y VDD LPPFET W=1.24U L=0.12U M=1 
X12 VDD C hnet19 VDD LPPFET W=1.24U L=0.12U M=1 
X13 hnet19 B hnet20 VDD LPPFET W=1.24U L=0.12U M=1 
X14 hnet20 A Y VDD LPPFET W=1.24U L=0.12U M=1 
X15 VDD C hnet9 VDD LPPFET W=1.24U L=0.12U M=1 
X16 hnet9 B hnet10 VDD LPPFET W=1.24U L=0.12U M=1 
X17 hnet10 A Y VDD LPPFET W=1.24U L=0.12U M=1 
X2 Y A VSS VSS LPNFET W=2.76U L=0.12U M=1 
X3 VDD C hnet21 VDD LPPFET W=1.24U L=0.12U M=1 
X4 hnet21 B hnet22 VDD LPPFET W=1.24U L=0.12U M=1 
X5 hnet22 A Y VDD LPPFET W=1.24U L=0.12U M=1 
X6 VDD C hnet11 VDD LPPFET W=1.24U L=0.12U M=1 
X7 hnet11 B hnet13 VDD LPPFET W=1.24U L=0.12U M=1 
X8 hnet13 A Y VDD LPPFET W=1.24U L=0.12U M=1 
X9 VDD C hnet7 VDD LPPFET W=1.24U L=0.12U M=1 
.ENDS NOR3X6TS 

**** 
*.SUBCKT NOR3X8TS Y A B C 
.SUBCKT NOR3X8TS Y A B C VSS VDD
X0 Y C VSS VSS LPNFET W=3.68U L=0.12U M=1 
X1 Y B VSS VSS LPNFET W=3.68U L=0.12U M=1 
X10 hnet7 B hnet19 VDD LPPFET W=1.28U L=0.12U M=1 
X11 hnet19 A Y VDD LPPFET W=1.28U L=0.12U M=1 
X12 VDD C hnet18 VDD LPPFET W=1.28U L=0.12U M=1 
X13 hnet18 B hnet12 VDD LPPFET W=1.28U L=0.12U M=1 
X14 hnet12 A Y VDD LPPFET W=1.28U L=0.12U M=1 
X15 VDD C hnet10 VDD LPPFET W=1.28U L=0.12U M=1 
X16 hnet10 B hnet8 VDD LPPFET W=1.28U L=0.12U M=1 
X17 hnet8 A Y VDD LPPFET W=1.28U L=0.12U M=1 
X18 VDD C hnet22 VDD LPPFET W=1.28U L=0.12U M=1 
X19 hnet22 B hnet21 VDD LPPFET W=1.28U L=0.12U M=1 
X2 Y A VSS VSS LPNFET W=3.68U L=0.12U M=1 
X20 hnet21 A Y VDD LPPFET W=1.28U L=0.12U M=1 
X3 VDD C hnet23 VDD LPPFET W=1.28U L=0.12U M=1 
X4 hnet23 B hnet24 VDD LPPFET W=1.28U L=0.12U M=1 
X5 hnet24 A Y VDD LPPFET W=1.28U L=0.12U M=1 
X6 VDD C hnet20 VDD LPPFET W=1.28U L=0.12U M=1 
X7 hnet20 B hnet9 VDD LPPFET W=1.28U L=0.12U M=1 
X8 hnet9 A Y VDD LPPFET W=1.28U L=0.12U M=1 
X9 VDD C hnet7 VDD LPPFET W=1.28U L=0.12U M=1 
.ENDS NOR3X8TS 

**** 
*.SUBCKT NOR3XLTS Y A B C 
.SUBCKT NOR3XLTS Y A B C VSS VDD
X0 Y C VSS VSS LPNFET W=0.24U L=0.12U M=1 
X1 Y B VSS VSS LPNFET W=0.24U L=0.12U M=1 
X2 Y A VSS VSS LPNFET W=0.24U L=0.12U M=1 
X3 VDD C hnet14 VDD LPPFET W=0.54U L=0.12U M=1 
X4 hnet14 B hnet13 VDD LPPFET W=0.54U L=0.12U M=1 
X5 hnet13 A Y VDD LPPFET W=0.54U L=0.12U M=1 
.ENDS NOR3XLTS 

**** 
*.SUBCKT NOR4BBX1TS Y AN BN C D 
.SUBCKT NOR4BBX1TS Y AN BN C D VSS VDD
X0 Y D VSS VSS LPNFET W=0.46U L=0.12U M=1 
X1 Y C VSS VSS LPNFET W=0.46U L=0.12U M=1 
X10 VDD AN nmin1 VDD LPPFET W=0.38U L=0.12U M=1 
X11 nmin1 AN VSS VSS LPNFET W=0.28U L=0.12U M=1 
X2 Y nmin2 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X3 Y nmin1 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X4 VDD D hnet13 VDD LPPFET W=1.2U L=0.12U M=1 
X5 hnet13 C hnet17 VDD LPPFET W=1.2U L=0.12U M=1 
X6 hnet17 nmin2 hnet11 VDD LPPFET W=1.2U L=0.12U M=1 
X7 hnet11 nmin1 Y VDD LPPFET W=1.2U L=0.12U M=1 
X8 VDD BN nmin2 VDD LPPFET W=0.38U L=0.12U M=1 
X9 nmin2 BN VSS VSS LPNFET W=0.28U L=0.12U M=1 
.ENDS NOR4BBX1TS 

**** 
*.SUBCKT NOR4BBX2TS Y AN BN C D 
.SUBCKT NOR4BBX2TS Y AN BN C D VSS VDD
X0 Y D VSS VSS LPNFET W=0.88U L=0.12U M=1 
X1 Y C VSS VSS LPNFET W=0.88U L=0.12U M=1 
X10 hnet10 nmin2 hnet21 VDD LPPFET W=1.04U L=0.12U M=1 
X11 hnet21 nmin1 Y VDD LPPFET W=1.04U L=0.12U M=1 
X12 VDD BN nmin2 VDD LPPFET W=0.78U L=0.12U M=1 
X13 nmin2 BN VSS VSS LPNFET W=0.56U L=0.12U M=1 
X14 VDD AN nmin1 VDD LPPFET W=0.78U L=0.12U M=1 
X15 nmin1 AN VSS VSS LPNFET W=0.56U L=0.12U M=1 
X2 Y nmin2 VSS VSS LPNFET W=0.88U L=0.12U M=1 
X3 Y nmin1 VSS VSS LPNFET W=0.88U L=0.12U M=1 
X4 VDD D hnet16 VDD LPPFET W=1.04U L=0.12U M=1 
X5 hnet16 C hnet15 VDD LPPFET W=1.04U L=0.12U M=1 
X6 hnet15 nmin2 hnet13 VDD LPPFET W=1.04U L=0.12U M=1 
X7 hnet13 nmin1 Y VDD LPPFET W=1.04U L=0.12U M=1 
X8 VDD D hnet11 VDD LPPFET W=1.04U L=0.12U M=1 
X9 hnet11 C hnet10 VDD LPPFET W=1.04U L=0.12U M=1 
.ENDS NOR4BBX2TS 

**** 
*.SUBCKT NOR4BBX4TS Y AN BN C D 
.SUBCKT NOR4BBX4TS Y AN BN C D VSS VDD
X0 Y D VSS VSS LPNFET W=1.68U L=0.12U M=1 
X1 Y C VSS VSS LPNFET W=1.68U L=0.12U M=1 
X10 hnet10 nmin2 hnet20 VDD LPPFET W=1.02U L=0.12U M=1 
X11 hnet20 nmin1 Y VDD LPPFET W=1.02U L=0.12U M=1 
X12 VDD D hnet18 VDD LPPFET W=1.02U L=0.12U M=1 
X13 hnet18 C hnet13 VDD LPPFET W=1.02U L=0.12U M=1 
X14 hnet13 nmin2 hnet15 VDD LPPFET W=1.02U L=0.12U M=1 
X15 hnet15 nmin1 Y VDD LPPFET W=1.02U L=0.12U M=1 
X16 VDD D hnet11 VDD LPPFET W=1.02U L=0.12U M=1 
X17 hnet11 C hnet26 VDD LPPFET W=1.02U L=0.12U M=1 
X18 hnet26 nmin2 hnet28 VDD LPPFET W=1.02U L=0.12U M=1 
X19 hnet28 nmin1 Y VDD LPPFET W=1.02U L=0.12U M=1 
X2 Y nmin2 VSS VSS LPNFET W=1.68U L=0.12U M=1 
X20 VDD BN nmin2 VDD LPPFET W=1.3U L=0.12U M=1 
X21 nmin2 BN VSS VSS LPNFET W=0.92U L=0.12U M=1 
X22 VDD AN nmin1 VDD LPPFET W=1.3U L=0.12U M=1 
X23 nmin1 AN VSS VSS LPNFET W=0.92U L=0.12U M=1 
X3 Y nmin1 VSS VSS LPNFET W=1.68U L=0.12U M=1 
X4 VDD D hnet17 VDD LPPFET W=1.02U L=0.12U M=1 
X5 hnet17 C hnet22 VDD LPPFET W=1.02U L=0.12U M=1 
X6 hnet22 nmin2 hnet21 VDD LPPFET W=1.02U L=0.12U M=1 
X7 hnet21 nmin1 Y VDD LPPFET W=1.02U L=0.12U M=1 
X8 VDD D hnet12 VDD LPPFET W=1.02U L=0.12U M=1 
X9 hnet12 C hnet10 VDD LPPFET W=1.02U L=0.12U M=1 
.ENDS NOR4BBX4TS 

**** 
*.SUBCKT NOR4BBXLTS Y AN BN C D 
.SUBCKT NOR4BBXLTS Y AN BN C D VSS VDD
X0 Y D VSS VSS LPNFET W=0.24U L=0.12U M=1 
X1 Y C VSS VSS LPNFET W=0.24U L=0.12U M=1 
X10 VDD AN nmin1 VDD LPPFET W=0.28U L=0.12U M=1 
X11 nmin1 AN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 Y nmin2 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X3 Y nmin1 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X4 VDD D hnet13 VDD LPPFET W=0.62U L=0.12U M=1 
X5 hnet13 C hnet17 VDD LPPFET W=0.62U L=0.12U M=1 
X6 hnet17 nmin2 hnet11 VDD LPPFET W=0.62U L=0.12U M=1 
X7 hnet11 nmin1 Y VDD LPPFET W=0.62U L=0.12U M=1 
X8 VDD BN nmin2 VDD LPPFET W=0.28U L=0.12U M=1 
X9 nmin2 BN VSS VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS NOR4BBXLTS 

**** 
*.SUBCKT NOR4BX1TS Y AN B C D 
.SUBCKT NOR4BX1TS Y AN B C D VSS VDD
X0 Y D VSS VSS LPNFET W=0.46U L=0.12U M=1 
X1 Y C VSS VSS LPNFET W=0.46U L=0.12U M=1 
X2 Y B VSS VSS LPNFET W=0.46U L=0.12U M=1 
X3 Y nmin1 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X4 VDD D hnet12 VDD LPPFET W=1.2U L=0.12U M=1 
X5 hnet12 C hnet16 VDD LPPFET W=1.2U L=0.12U M=1 
X6 hnet16 B hnet10 VDD LPPFET W=1.2U L=0.12U M=1 
X7 hnet10 nmin1 Y VDD LPPFET W=1.2U L=0.12U M=1 
X8 VDD AN nmin1 VDD LPPFET W=0.38U L=0.12U M=1 
X9 nmin1 AN VSS VSS LPNFET W=0.28U L=0.12U M=1 
.ENDS NOR4BX1TS 

**** 
*.SUBCKT NOR4BX2TS Y AN B C D 
.SUBCKT NOR4BX2TS Y AN B C D VSS VDD
X0 Y D VSS VSS LPNFET W=0.92U L=0.12U M=1 
X1 Y C VSS VSS LPNFET W=0.92U L=0.12U M=1 
X10 hnet9 B hnet20 VDD LPPFET W=1.12U L=0.12U M=1 
X11 hnet20 nmin1 Y VDD LPPFET W=1.12U L=0.12U M=1 
X12 VDD AN nmin1 VDD LPPFET W=0.78U L=0.12U M=1 
X13 nmin1 AN VSS VSS LPNFET W=0.56U L=0.12U M=1 
X2 Y B VSS VSS LPNFET W=0.92U L=0.12U M=1 
X3 Y nmin1 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X4 VDD D hnet15 VDD LPPFET W=1.12U L=0.12U M=1 
X5 hnet15 C hnet14 VDD LPPFET W=1.12U L=0.12U M=1 
X6 hnet14 B hnet12 VDD LPPFET W=1.12U L=0.12U M=1 
X7 hnet12 nmin1 Y VDD LPPFET W=1.12U L=0.12U M=1 
X8 VDD D hnet10 VDD LPPFET W=1.12U L=0.12U M=1 
X9 hnet10 C hnet9 VDD LPPFET W=1.12U L=0.12U M=1 
.ENDS NOR4BX2TS 

**** 
*.SUBCKT NOR4BX4TS Y AN B C D 
.SUBCKT NOR4BX4TS Y AN B C D VSS VDD
X0 Y D VSS VSS LPNFET W=1.68U L=0.12U M=1 
X1 Y C VSS VSS LPNFET W=1.68U L=0.12U M=1 
X10 hnet9 B hnet19 VDD LPPFET W=1.02U L=0.12U M=1 
X11 hnet19 nmin1 Y VDD LPPFET W=1.02U L=0.12U M=1 
X12 VDD D hnet17 VDD LPPFET W=1.02U L=0.12U M=1 
X13 hnet17 C hnet12 VDD LPPFET W=1.02U L=0.12U M=1 
X14 hnet12 B hnet14 VDD LPPFET W=1.02U L=0.12U M=1 
X15 hnet14 nmin1 Y VDD LPPFET W=1.02U L=0.12U M=1 
X16 VDD D hnet10 VDD LPPFET W=1.02U L=0.12U M=1 
X17 hnet10 C hnet25 VDD LPPFET W=1.02U L=0.12U M=1 
X18 hnet25 B hnet27 VDD LPPFET W=1.02U L=0.12U M=1 
X19 hnet27 nmin1 Y VDD LPPFET W=1.02U L=0.12U M=1 
X2 Y B VSS VSS LPNFET W=1.68U L=0.12U M=1 
X20 VDD AN nmin1 VDD LPPFET W=1.3U L=0.12U M=1 
X21 nmin1 AN VSS VSS LPNFET W=0.92U L=0.12U M=1 
X3 Y nmin1 VSS VSS LPNFET W=1.68U L=0.12U M=1 
X4 VDD D hnet16 VDD LPPFET W=1.02U L=0.12U M=1 
X5 hnet16 C hnet21 VDD LPPFET W=1.02U L=0.12U M=1 
X6 hnet21 B hnet20 VDD LPPFET W=1.02U L=0.12U M=1 
X7 hnet20 nmin1 Y VDD LPPFET W=1.02U L=0.12U M=1 
X8 VDD D hnet11 VDD LPPFET W=1.02U L=0.12U M=1 
X9 hnet11 C hnet9 VDD LPPFET W=1.02U L=0.12U M=1 
.ENDS NOR4BX4TS 

**** 
*.SUBCKT NOR4BXLTS Y AN B C D 
.SUBCKT NOR4BXLTS Y AN B C D VSS VDD
X0 Y D VSS VSS LPNFET W=0.24U L=0.12U M=1 
X1 Y C VSS VSS LPNFET W=0.24U L=0.12U M=1 
X2 Y B VSS VSS LPNFET W=0.24U L=0.12U M=1 
X3 Y nmin1 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X4 VDD D hnet12 VDD LPPFET W=0.62U L=0.12U M=1 
X5 hnet12 C hnet16 VDD LPPFET W=0.62U L=0.12U M=1 
X6 hnet16 B hnet10 VDD LPPFET W=0.62U L=0.12U M=1 
X7 hnet10 nmin1 Y VDD LPPFET W=0.62U L=0.12U M=1 
X8 VDD AN nmin1 VDD LPPFET W=0.28U L=0.12U M=1 
X9 nmin1 AN VSS VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS NOR4BXLTS 

**** 
*.SUBCKT NOR4X1TS Y A B C D 
.SUBCKT NOR4X1TS Y A B C D VSS VDD
X0 Y D VSS VSS LPNFET W=0.46U L=0.12U M=1 
X1 Y C VSS VSS LPNFET W=0.46U L=0.12U M=1 
X2 Y B VSS VSS LPNFET W=0.46U L=0.12U M=1 
X3 Y A VSS VSS LPNFET W=0.46U L=0.12U M=1 
X4 VDD D hnet11 VDD LPPFET W=1.2U L=0.12U M=1 
X5 hnet11 C hnet15 VDD LPPFET W=1.2U L=0.12U M=1 
X6 hnet15 B hnet9 VDD LPPFET W=1.2U L=0.12U M=1 
X7 hnet9 A Y VDD LPPFET W=1.2U L=0.12U M=1 
.ENDS NOR4X1TS 

**** 
*.SUBCKT NOR4X2TS Y A B C D 
.SUBCKT NOR4X2TS Y A B C D VSS VDD
X0 Y D VSS VSS LPNFET W=0.92U L=0.12U M=1 
X1 Y C VSS VSS LPNFET W=0.92U L=0.12U M=1 
X10 hnet8 B hnet19 VDD LPPFET W=1.2U L=0.12U M=1 
X11 hnet19 A Y VDD LPPFET W=1.2U L=0.12U M=1 
X2 Y B VSS VSS LPNFET W=0.92U L=0.12U M=1 
X3 Y A VSS VSS LPNFET W=0.92U L=0.12U M=1 
X4 VDD D hnet14 VDD LPPFET W=1.2U L=0.12U M=1 
X5 hnet14 C hnet13 VDD LPPFET W=1.2U L=0.12U M=1 
X6 hnet13 B hnet11 VDD LPPFET W=1.2U L=0.12U M=1 
X7 hnet11 A Y VDD LPPFET W=1.2U L=0.12U M=1 
X8 VDD D hnet9 VDD LPPFET W=1.2U L=0.12U M=1 
X9 hnet9 C hnet8 VDD LPPFET W=1.2U L=0.12U M=1 
.ENDS NOR4X2TS 

**** 
*.SUBCKT NOR4X4TS Y A B C D 
.SUBCKT NOR4X4TS Y A B C D VSS VDD
X0 Y D VSS VSS LPNFET W=1.68U L=0.12U M=1 
X1 Y C VSS VSS LPNFET W=1.68U L=0.12U M=1 
X10 hnet8 B hnet18 VDD LPPFET W=1.08U L=0.12U M=1 
X11 hnet18 A Y VDD LPPFET W=1.08U L=0.12U M=1 
X12 VDD D hnet16 VDD LPPFET W=1.08U L=0.12U M=1 
X13 hnet16 C hnet11 VDD LPPFET W=1.08U L=0.12U M=1 
X14 hnet11 B hnet13 VDD LPPFET W=1.08U L=0.12U M=1 
X15 hnet13 A Y VDD LPPFET W=1.08U L=0.12U M=1 
X16 VDD D hnet9 VDD LPPFET W=1.08U L=0.12U M=1 
X17 hnet9 C hnet24 VDD LPPFET W=1.08U L=0.12U M=1 
X18 hnet24 B hnet26 VDD LPPFET W=1.08U L=0.12U M=1 
X19 hnet26 A Y VDD LPPFET W=1.08U L=0.12U M=1 
X2 Y B VSS VSS LPNFET W=1.68U L=0.12U M=1 
X3 Y A VSS VSS LPNFET W=1.68U L=0.12U M=1 
X4 VDD D hnet15 VDD LPPFET W=1.08U L=0.12U M=1 
X5 hnet15 C hnet20 VDD LPPFET W=1.08U L=0.12U M=1 
X6 hnet20 B hnet19 VDD LPPFET W=1.08U L=0.12U M=1 
X7 hnet19 A Y VDD LPPFET W=1.08U L=0.12U M=1 
X8 VDD D hnet10 VDD LPPFET W=1.08U L=0.12U M=1 
X9 hnet10 C hnet8 VDD LPPFET W=1.08U L=0.12U M=1 
.ENDS NOR4X4TS 

**** 
*.SUBCKT NOR4X6TS Y A B C D 
.SUBCKT NOR4X6TS Y A B C D VSS VDD
X0 Y D VSS VSS LPNFET W=2.5U L=0.12U M=1 
X1 Y C VSS VSS LPNFET W=2.5U L=0.12U M=1 
X10 hnet8 B hnet12 VDD LPPFET W=1.04U L=0.12U M=1 
X11 hnet12 A Y VDD LPPFET W=1.04U L=0.12U M=1 
X12 VDD D hnet28 VDD LPPFET W=1.04U L=0.12U M=1 
X13 hnet28 C hnet27 VDD LPPFET W=1.04U L=0.12U M=1 
X14 hnet27 B hnet13 VDD LPPFET W=1.04U L=0.12U M=1 
X15 hnet13 A Y VDD LPPFET W=1.04U L=0.12U M=1 
X16 VDD D hnet10 VDD LPPFET W=1.04U L=0.12U M=1 
X17 hnet10 C hnet11 VDD LPPFET W=1.04U L=0.12U M=1 
X18 hnet11 B hnet32 VDD LPPFET W=1.04U L=0.12U M=1 
X19 hnet32 A Y VDD LPPFET W=1.04U L=0.12U M=1 
X2 Y B VSS VSS LPNFET W=2.5U L=0.12U M=1 
X20 VDD D hnet18 VDD LPPFET W=1.04U L=0.12U M=1 
X21 hnet18 C hnet19 VDD LPPFET W=1.04U L=0.12U M=1 
X22 hnet19 B hnet15 VDD LPPFET W=1.04U L=0.12U M=1 
X23 hnet15 A Y VDD LPPFET W=1.04U L=0.12U M=1 
X24 VDD D hnet30 VDD LPPFET W=1.04U L=0.12U M=1 
X25 hnet30 C hnet9 VDD LPPFET W=1.04U L=0.12U M=1 
X26 hnet9 B hnet23 VDD LPPFET W=1.04U L=0.12U M=1 
X27 hnet23 A Y VDD LPPFET W=1.04U L=0.12U M=1 
X3 Y A VSS VSS LPNFET W=2.5U L=0.12U M=1 
X4 VDD D hnet31 VDD LPPFET W=1.04U L=0.12U M=1 
X5 hnet31 C hnet21 VDD LPPFET W=1.04U L=0.12U M=1 
X6 hnet21 B hnet17 VDD LPPFET W=1.04U L=0.12U M=1 
X7 hnet17 A Y VDD LPPFET W=1.04U L=0.12U M=1 
X8 VDD D hnet14 VDD LPPFET W=1.04U L=0.12U M=1 
X9 hnet14 C hnet8 VDD LPPFET W=1.04U L=0.12U M=1 
.ENDS NOR4X6TS 

**** 
*.SUBCKT NOR4X8TS Y A B C D 
.SUBCKT NOR4X8TS Y A B C D VSS VDD
X0 Y D VSS VSS LPNFET W=3.36U L=0.12U M=1 
X1 Y C VSS VSS LPNFET W=3.36U L=0.12U M=1 
X10 hnet17 B hnet12 VDD LPPFET W=1.04U L=0.12U M=1 
X11 hnet12 A Y VDD LPPFET W=1.04U L=0.12U M=1 
X12 VDD D hnet34 VDD LPPFET W=1.04U L=0.12U M=1 
X13 hnet34 C hnet36 VDD LPPFET W=1.04U L=0.12U M=1 
X14 hnet36 B hnet15 VDD LPPFET W=1.04U L=0.12U M=1 
X15 hnet15 A Y VDD LPPFET W=1.04U L=0.12U M=1 
X16 VDD D hnet11 VDD LPPFET W=1.04U L=0.12U M=1 
X17 hnet11 C hnet37 VDD LPPFET W=1.04U L=0.12U M=1 
X18 hnet37 B hnet8 VDD LPPFET W=1.04U L=0.12U M=1 
X19 hnet8 A Y VDD LPPFET W=1.04U L=0.12U M=1 
X2 Y B VSS VSS LPNFET W=3.36U L=0.12U M=1 
X20 VDD D hnet19 VDD LPPFET W=1.04U L=0.12U M=1 
X21 hnet19 C hnet16 VDD LPPFET W=1.04U L=0.12U M=1 
X22 hnet16 B hnet20 VDD LPPFET W=1.04U L=0.12U M=1 
X23 hnet20 A Y VDD LPPFET W=1.04U L=0.12U M=1 
X24 VDD D hnet13 VDD LPPFET W=1.04U L=0.12U M=1 
X25 hnet13 C hnet10 VDD LPPFET W=1.04U L=0.12U M=1 
X26 hnet10 B hnet27 VDD LPPFET W=1.04U L=0.12U M=1 
X27 hnet27 A Y VDD LPPFET W=1.04U L=0.12U M=1 
X28 VDD D hnet25 VDD LPPFET W=1.04U L=0.12U M=1 
X29 hnet25 C hnet23 VDD LPPFET W=1.04U L=0.12U M=1 
X3 Y A VSS VSS LPNFET W=3.36U L=0.12U M=1 
X30 hnet23 B hnet22 VDD LPPFET W=1.04U L=0.12U M=1 
X31 hnet22 A Y VDD LPPFET W=1.04U L=0.12U M=1 
X32 VDD D hnet33 VDD LPPFET W=1.04U L=0.12U M=1 
X33 hnet33 C hnet21 VDD LPPFET W=1.04U L=0.12U M=1 
X34 hnet21 B hnet14 VDD LPPFET W=1.04U L=0.12U M=1 
X35 hnet14 A Y VDD LPPFET W=1.04U L=0.12U M=1 
X4 VDD D hnet29 VDD LPPFET W=1.04U L=0.12U M=1 
X5 hnet29 C hnet35 VDD LPPFET W=1.04U L=0.12U M=1 
X6 hnet35 B hnet26 VDD LPPFET W=1.04U L=0.12U M=1 
X7 hnet26 A Y VDD LPPFET W=1.04U L=0.12U M=1 
X8 VDD D hnet9 VDD LPPFET W=1.04U L=0.12U M=1 
X9 hnet9 C hnet17 VDD LPPFET W=1.04U L=0.12U M=1 
.ENDS NOR4X8TS 

**** 
*.SUBCKT NOR4XLTS Y A B C D 
.SUBCKT NOR4XLTS Y A B C D VSS VDD
X0 Y D VSS VSS LPNFET W=0.24U L=0.12U M=1 
X1 Y C VSS VSS LPNFET W=0.24U L=0.12U M=1 
X2 Y B VSS VSS LPNFET W=0.24U L=0.12U M=1 
X3 Y A VSS VSS LPNFET W=0.24U L=0.12U M=1 
X4 VDD D hnet11 VDD LPPFET W=0.62U L=0.12U M=1 
X5 hnet11 C hnet15 VDD LPPFET W=0.62U L=0.12U M=1 
X6 hnet15 B hnet9 VDD LPPFET W=0.62U L=0.12U M=1 
X7 hnet9 A Y VDD LPPFET W=0.62U L=0.12U M=1 
.ENDS NOR4XLTS 

**** 
*.SUBCKT OA21X1TS Y A0 A1 B0 
.SUBCKT OA21X1TS Y A0 A1 B0 VSS VDD
X0 VDD nmin Y VDD LPPFET W=0.64U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=0.46U L=0.12U M=1 
X2 VDD A1 hnet16 VDD LPPFET W=0.34U L=0.12U M=1 
X3 hnet16 A0 nmin VDD LPPFET W=0.34U L=0.12U M=1 
X4 nmin B0 net27 VSS LPNFET W=0.26U L=0.12U M=1 
X5 net27 A1 VSS VSS LPNFET W=0.26U L=0.12U M=1 
X6 net27 A0 VSS VSS LPNFET W=0.26U L=0.12U M=1 
X7 nmin B0 VDD VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS OA21X1TS 

**** 
*.SUBCKT OA21X2TS Y A0 A1 B0 
.SUBCKT OA21X2TS Y A0 A1 B0 VSS VDD
X0 VDD nmin Y VDD LPPFET W=1.28U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=0.92U L=0.12U M=1 
X2 VDD A1 hnet16 VDD LPPFET W=0.68U L=0.12U M=1 
X3 hnet16 A0 nmin VDD LPPFET W=0.68U L=0.12U M=1 
X4 nmin B0 net27 VSS LPNFET W=0.5U L=0.12U M=1 
X5 net27 A1 VSS VSS LPNFET W=0.5U L=0.12U M=1 
X6 net27 A0 VSS VSS LPNFET W=0.5U L=0.12U M=1 
X7 nmin B0 VDD VDD LPPFET W=0.52U L=0.12U M=1 
.ENDS OA21X2TS 

**** 
*.SUBCKT OA21X4TS Y A0 A1 B0 
.SUBCKT OA21X4TS Y A0 A1 B0 VSS VDD
X0 VDD nmin Y VDD LPPFET W=2.58U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=1.7U L=0.12U M=1 
X2 VDD A1 hnet16 VDD LPPFET W=1.3U L=0.12U M=1 
X3 hnet16 A0 nmin VDD LPPFET W=1.3U L=0.12U M=1 
X4 nmin B0 net27 VSS LPNFET W=0.92U L=0.12U M=1 
X5 net27 A1 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X6 net27 A0 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X7 nmin B0 VDD VDD LPPFET W=1.02U L=0.12U M=1 
.ENDS OA21X4TS 

**** 
*.SUBCKT OA21XLTS Y A0 A1 B0 
.SUBCKT OA21XLTS Y A0 A1 B0 VSS VDD
X0 VDD nmin Y VDD LPPFET W=0.42U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=0.24U L=0.12U M=1 
X2 VDD A1 hnet16 VDD LPPFET W=0.3U L=0.12U M=1 
X3 hnet16 A0 nmin VDD LPPFET W=0.3U L=0.12U M=1 
X4 nmin B0 net27 VSS LPNFET W=0.26U L=0.12U M=1 
X5 net27 A1 VSS VSS LPNFET W=0.26U L=0.12U M=1 
X6 net27 A0 VSS VSS LPNFET W=0.26U L=0.12U M=1 
X7 nmin B0 VDD VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS OA21XLTS 

**** 
*.SUBCKT OA22X1TS Y A0 A1 B0 B1 
.SUBCKT OA22X1TS Y A0 A1 B0 B1 VSS VDD
X0 VDD nmin Y VDD LPPFET W=0.64U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=0.46U L=0.12U M=1 
X2 VDD B1 hnet17 VDD LPPFET W=0.34U L=0.12U M=1 
X3 hnet17 B0 nmin VDD LPPFET W=0.34U L=0.12U M=1 
X4 VDD A1 hnet21 VDD LPPFET W=0.34U L=0.12U M=1 
X5 hnet21 A0 nmin VDD LPPFET W=0.34U L=0.12U M=1 
X6 nmin A0 net40 VSS LPNFET W=0.24U L=0.12U M=1 
X7 nmin A1 net40 VSS LPNFET W=0.24U L=0.12U M=1 
X8 net40 B0 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X9 net40 B1 VSS VSS LPNFET W=0.24U L=0.12U M=1 
.ENDS OA22X1TS 

**** 
*.SUBCKT OA22X2TS Y A0 A1 B0 B1 
.SUBCKT OA22X2TS Y A0 A1 B0 B1 VSS VDD
X0 VDD nmin Y VDD LPPFET W=1.28U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=0.92U L=0.12U M=1 
X2 VDD B1 hnet17 VDD LPPFET W=0.68U L=0.12U M=1 
X3 hnet17 B0 nmin VDD LPPFET W=0.68U L=0.12U M=1 
X4 VDD A1 hnet21 VDD LPPFET W=0.68U L=0.12U M=1 
X5 hnet21 A0 nmin VDD LPPFET W=0.68U L=0.12U M=1 
X6 nmin A0 net40 VSS LPNFET W=0.48U L=0.12U M=1 
X7 nmin A1 net40 VSS LPNFET W=0.48U L=0.12U M=1 
X8 net40 B0 VSS VSS LPNFET W=0.48U L=0.12U M=1 
X9 net40 B1 VSS VSS LPNFET W=0.48U L=0.12U M=1 
.ENDS OA22X2TS 

**** 
*.SUBCKT OA22X4TS Y A0 A1 B0 B1 
.SUBCKT OA22X4TS Y A0 A1 B0 B1 VSS VDD
X0 VDD nmin Y VDD LPPFET W=2.4U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=1.84U L=0.12U M=1 
X2 VDD B1 hnet17 VDD LPPFET W=1.2U L=0.12U M=1 
X3 hnet17 B0 nmin VDD LPPFET W=1.2U L=0.12U M=1 
X4 VDD A1 hnet21 VDD LPPFET W=1.2U L=0.12U M=1 
X5 hnet21 A0 nmin VDD LPPFET W=1.2U L=0.12U M=1 
X6 nmin A0 net40 VSS LPNFET W=0.92U L=0.12U M=1 
X7 nmin A1 net40 VSS LPNFET W=0.92U L=0.12U M=1 
X8 net40 B0 VSS VSS LPNFET W=0.78U L=0.12U M=1 
X9 net40 B1 VSS VSS LPNFET W=0.92U L=0.12U M=1 
.ENDS OA22X4TS 

**** 
*.SUBCKT OA22XLTS Y A0 A1 B0 B1 
.SUBCKT OA22XLTS Y A0 A1 B0 B1 VSS VDD
X0 VDD nmin Y VDD LPPFET W=0.42U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=0.24U L=0.12U M=1 
X2 VDD B1 hnet17 VDD LPPFET W=0.3U L=0.12U M=1 
X3 hnet17 B0 nmin VDD LPPFET W=0.3U L=0.12U M=1 
X4 VDD A1 hnet21 VDD LPPFET W=0.3U L=0.12U M=1 
X5 hnet21 A0 nmin VDD LPPFET W=0.3U L=0.12U M=1 
X6 nmin A0 net40 VSS LPNFET W=0.26U L=0.12U M=1 
X7 nmin A1 net40 VSS LPNFET W=0.26U L=0.12U M=1 
X8 net40 B0 VSS VSS LPNFET W=0.26U L=0.12U M=1 
X9 net40 B1 VSS VSS LPNFET W=0.26U L=0.12U M=1 
.ENDS OA22XLTS 

**** 
*.SUBCKT OAI211X1TS Y A0 A1 B0 C0 
.SUBCKT OAI211X1TS Y A0 A1 B0 C0 VSS VDD
X0 VDD A1 hnet15 VDD LPPFET W=0.84U L=0.12U M=1 
X1 hnet15 A0 Y VDD LPPFET W=0.84U L=0.12U M=1 
X2 net25 C0 net32 VSS LPNFET W=0.72U L=0.12U M=1 
X3 Y B0 net25 VSS LPNFET W=0.72U L=0.12U M=1 
X4 net32 A1 VSS VSS LPNFET W=0.72U L=0.12U M=1 
X5 net32 A0 VSS VSS LPNFET W=0.72U L=0.12U M=1 
X6 Y C0 VDD VDD LPPFET W=0.64U L=0.12U M=1 
X7 Y B0 VDD VDD LPPFET W=0.64U L=0.12U M=1 
.ENDS OAI211X1TS 

**** 
*.SUBCKT OAI211X2TS Y A0 A1 B0 C0 
.SUBCKT OAI211X2TS Y A0 A1 B0 C0 VSS VDD
X0 VDD A1 hnet17 VDD LPPFET W=0.84U L=0.12U M=1 
X1 hnet17 A0 Y VDD LPPFET W=0.84U L=0.12U M=1 
X10 Y C0 VDD VDD LPPFET W=1.28U L=0.12U M=1 
X11 Y B0 VDD VDD LPPFET W=1.28U L=0.12U M=1 
X2 VDD A1 hnet14 VDD LPPFET W=0.84U L=0.12U M=1 
X3 hnet14 A0 Y VDD LPPFET W=0.84U L=0.12U M=1 
X4 net25 C0 net38 VSS LPNFET W=0.58U L=0.12U M=1 
X5 Y B0 net25 VSS LPNFET W=0.58U L=0.12U M=1 
X6 net31 C0 net38 VSS LPNFET W=0.58U L=0.12U M=1 
X7 Y B0 net31 VSS LPNFET W=0.58U L=0.12U M=1 
X8 net38 A1 VSS VSS LPNFET W=1.32U L=0.12U M=1 
X9 net38 A0 VSS VSS LPNFET W=1.32U L=0.12U M=1 
.ENDS OAI211X2TS 

**** 
*.SUBCKT OAI211X4TS Y A0 A1 B0 C0 
.SUBCKT OAI211X4TS Y A0 A1 B0 C0 VSS VDD
X0 VDD net23 net19 VDD LPPFET W=1.02U L=0.12U M=1 
X1 net19 net23 VSS VSS LPNFET W=0.74U L=0.12U M=1 
X10 net23 C0 VDD VDD LPPFET W=0.4U L=0.12U M=1 
X11 net23 B0 VDD VDD LPPFET W=0.4U L=0.12U M=1 
X2 VDD net19 Y VDD LPPFET W=2.56U L=0.12U M=1 
X3 Y net19 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X4 VDD A1 hnet21 VDD LPPFET W=0.54U L=0.12U M=1 
X5 hnet21 A0 net23 VDD LPPFET W=0.54U L=0.12U M=1 
X6 net30 C0 net37 VSS LPNFET W=0.46U L=0.12U M=1 
X7 net23 B0 net30 VSS LPNFET W=0.46U L=0.12U M=1 
X8 net37 A1 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X9 net37 A0 VSS VSS LPNFET W=0.46U L=0.12U M=1 
.ENDS OAI211X4TS 

**** 
*.SUBCKT OAI211XLTS Y A0 A1 B0 C0 
.SUBCKT OAI211XLTS Y A0 A1 B0 C0 VSS VDD
X0 VDD A1 hnet15 VDD LPPFET W=0.44U L=0.12U M=1 
X1 hnet15 A0 Y VDD LPPFET W=0.44U L=0.12U M=1 
X2 net25 C0 net32 VSS LPNFET W=0.48U L=0.12U M=1 
X3 Y B0 net25 VSS LPNFET W=0.48U L=0.12U M=1 
X4 net32 A1 VSS VSS LPNFET W=0.48U L=0.12U M=1 
X5 net32 A0 VSS VSS LPNFET W=0.48U L=0.12U M=1 
X6 Y C0 VDD VDD LPPFET W=0.42U L=0.12U M=1 
X7 Y B0 VDD VDD LPPFET W=0.42U L=0.12U M=1 
.ENDS OAI211XLTS 

**** 
*.SUBCKT OAI21X1TS Y A0 A1 B0 
.SUBCKT OAI21X1TS Y A0 A1 B0 VSS VDD
X0 VDD A1 hnet13 VDD LPPFET W=0.84U L=0.12U M=1 
X1 hnet13 A0 Y VDD LPPFET W=0.84U L=0.12U M=1 
X2 Y B0 net25 VSS LPNFET W=0.6U L=0.12U M=1 
X3 net25 A1 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X4 net25 A0 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X5 Y B0 VDD VDD LPPFET W=0.64U L=0.12U M=1 
.ENDS OAI21X1TS 

**** 
*.SUBCKT OAI21X2TS Y A0 A1 B0 
.SUBCKT OAI21X2TS Y A0 A1 B0 VSS VDD
X0 VDD A1 hnet14 VDD LPPFET W=0.84U L=0.12U M=1 
X1 hnet14 A0 Y VDD LPPFET W=0.84U L=0.12U M=1 
X2 VDD A1 hnet11 VDD LPPFET W=0.84U L=0.12U M=1 
X3 hnet11 A0 Y VDD LPPFET W=0.84U L=0.12U M=1 
X4 Y B0 net25 VSS LPNFET W=1.22U L=0.12U M=1 
X5 net25 A1 VSS VSS LPNFET W=1.22U L=0.12U M=1 
X6 net25 A0 VSS VSS LPNFET W=1.22U L=0.12U M=1 
X7 Y B0 VDD VDD LPPFET W=1.28U L=0.12U M=1 
.ENDS OAI21X2TS 

**** 
*.SUBCKT OAI21X4TS Y A0 A1 B0 
.SUBCKT OAI21X4TS Y A0 A1 B0 VSS VDD
X0 VDD A1 hnet14 VDD LPPFET W=1.12U L=0.12U M=1 
X1 hnet14 A0 Y VDD LPPFET W=1.12U L=0.12U M=1 
X2 VDD A1 hnet11 VDD LPPFET W=1.12U L=0.12U M=1 
X3 hnet11 A0 Y VDD LPPFET W=1.12U L=0.12U M=1 
X4 VDD A1 hnet10 VDD LPPFET W=1.12U L=0.12U M=1 
X5 hnet10 A0 Y VDD LPPFET W=1.12U L=0.12U M=1 
X6 Y B0 net25 VSS LPNFET W=2.46U L=0.12U M=1 
X7 net25 A1 VSS VSS LPNFET W=2.24U L=0.12U M=1 
X8 net25 A0 VSS VSS LPNFET W=2.24U L=0.12U M=1 
X9 Y B0 VDD VDD LPPFET W=2.56U L=0.12U M=1 
.ENDS OAI21X4TS 

**** 
*.SUBCKT OAI21XLTS Y A0 A1 B0 
.SUBCKT OAI21XLTS Y A0 A1 B0 VSS VDD
X0 VDD A1 hnet13 VDD LPPFET W=0.44U L=0.12U M=1 
X1 hnet13 A0 Y VDD LPPFET W=0.44U L=0.12U M=1 
X2 Y B0 net25 VSS LPNFET W=0.4U L=0.12U M=1 
X3 net25 A1 VSS VSS LPNFET W=0.4U L=0.12U M=1 
X4 net25 A0 VSS VSS LPNFET W=0.4U L=0.12U M=1 
X5 Y B0 VDD VDD LPPFET W=0.42U L=0.12U M=1 
.ENDS OAI21XLTS 

**** 
*.SUBCKT OAI221X1TS Y A0 A1 B0 B1 C0 
.SUBCKT OAI221X1TS Y A0 A1 B0 B1 C0 VSS VDD
X0 VDD B1 hnet16 VDD LPPFET W=0.84U L=0.12U M=1 
X1 hnet16 B0 Y VDD LPPFET W=0.84U L=0.12U M=1 
X2 VDD A1 hnet20 VDD LPPFET W=0.84U L=0.12U M=1 
X3 hnet20 A0 Y VDD LPPFET W=0.84U L=0.12U M=1 
X4 Y C0 VDD VDD LPPFET W=0.64U L=0.12U M=1 
X5 Y C0 net42 VSS LPNFET W=0.66U L=0.12U M=1 
X6 net42 A0 net48 VSS LPNFET W=0.66U L=0.12U M=1 
X7 net42 A1 net48 VSS LPNFET W=0.66U L=0.12U M=1 
X8 net48 B0 VSS VSS LPNFET W=0.72U L=0.12U M=1 
X9 net48 B1 VSS VSS LPNFET W=0.72U L=0.12U M=1 
.ENDS OAI221X1TS 

**** 
*.SUBCKT OAI221X2TS Y A0 A1 B0 B1 C0 
.SUBCKT OAI221X2TS Y A0 A1 B0 B1 C0 VSS VDD
X0 VDD B1 hnet17 VDD LPPFET W=0.84U L=0.12U M=1 
X1 hnet17 B0 Y VDD LPPFET W=0.84U L=0.12U M=1 
X10 net42 A0 net48 VSS LPNFET W=1.46U L=0.12U M=1 
X11 net42 A1 net48 VSS LPNFET W=1.46U L=0.12U M=1 
X12 net48 B0 VSS VSS LPNFET W=1.46U L=0.12U M=1 
X13 net48 B1 VSS VSS LPNFET W=1.46U L=0.12U M=1 
X2 VDD B1 hnet14 VDD LPPFET W=0.84U L=0.12U M=1 
X3 hnet14 B0 Y VDD LPPFET W=0.84U L=0.12U M=1 
X4 VDD A1 hnet22 VDD LPPFET W=0.76U L=0.12U M=1 
X5 hnet22 A0 Y VDD LPPFET W=0.76U L=0.12U M=1 
X6 VDD A1 hnet19 VDD LPPFET W=0.76U L=0.12U M=1 
X7 hnet19 A0 Y VDD LPPFET W=0.76U L=0.12U M=1 
X8 Y C0 VDD VDD LPPFET W=1.28U L=0.12U M=1 
X9 Y C0 net42 VSS LPNFET W=1.32U L=0.12U M=1 
.ENDS OAI221X2TS 

**** 
*.SUBCKT OAI221X4TS Y A0 A1 B0 B1 C0 
.SUBCKT OAI221X4TS Y A0 A1 B0 B1 C0 VSS VDD
X0 VDD net30 net26 VDD LPPFET W=1.02U L=0.12U M=1 
X1 net26 net30 VSS VSS LPNFET W=0.74U L=0.12U M=1 
X10 net47 A0 net53 VSS LPNFET W=0.46U L=0.12U M=1 
X11 net47 A1 net53 VSS LPNFET W=0.46U L=0.12U M=1 
X12 net53 B0 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X13 net53 B1 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X2 VDD net26 Y VDD LPPFET W=2.56U L=0.12U M=1 
X3 Y net26 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X4 VDD B1 hnet22 VDD LPPFET W=0.54U L=0.12U M=1 
X5 hnet22 B0 net30 VDD LPPFET W=0.54U L=0.12U M=1 
X6 VDD A1 hnet26 VDD LPPFET W=0.54U L=0.12U M=1 
X7 hnet26 A0 net30 VDD LPPFET W=0.54U L=0.12U M=1 
X8 net30 C0 VDD VDD LPPFET W=0.4U L=0.12U M=1 
X9 net30 C0 net47 VSS LPNFET W=0.44U L=0.12U M=1 
.ENDS OAI221X4TS 

**** 
*.SUBCKT OAI221XLTS Y A0 A1 B0 B1 C0 
.SUBCKT OAI221XLTS Y A0 A1 B0 B1 C0 VSS VDD
X0 VDD B1 hnet16 VDD LPPFET W=0.44U L=0.12U M=1 
X1 hnet16 B0 Y VDD LPPFET W=0.44U L=0.12U M=1 
X2 VDD A1 hnet20 VDD LPPFET W=0.44U L=0.12U M=1 
X3 hnet20 A0 Y VDD LPPFET W=0.44U L=0.12U M=1 
X4 Y C0 VDD VDD LPPFET W=0.42U L=0.12U M=1 
X5 Y C0 net42 VSS LPNFET W=0.48U L=0.12U M=1 
X6 net42 A0 net48 VSS LPNFET W=0.48U L=0.12U M=1 
X7 net42 A1 net48 VSS LPNFET W=0.48U L=0.12U M=1 
X8 net48 B0 VSS VSS LPNFET W=0.48U L=0.12U M=1 
X9 net48 B1 VSS VSS LPNFET W=0.48U L=0.12U M=1 
.ENDS OAI221XLTS 

**** 
*.SUBCKT OAI222X1TS Y A0 A1 B0 B1 C0 C1 
.SUBCKT OAI222X1TS Y A0 A1 B0 B1 C0 C1 VSS VDD
X0 VDD B1 hnet17 VDD LPPFET W=0.84U L=0.12U M=1 
X1 hnet17 B0 Y VDD LPPFET W=0.84U L=0.12U M=1 
X10 net55 B0 VSS VSS LPNFET W=0.66U L=0.12U M=1 
X11 net55 B1 VSS VSS LPNFET W=0.66U L=0.12U M=1 
X2 VDD A1 hnet22 VDD LPPFET W=0.84U L=0.12U M=1 
X3 hnet22 A0 Y VDD LPPFET W=0.84U L=0.12U M=1 
X4 VDD C1 hnet27 VDD LPPFET W=0.84U L=0.12U M=1 
X5 hnet27 C0 Y VDD LPPFET W=0.84U L=0.12U M=1 
X6 Y C0 net49 VSS LPNFET W=0.66U L=0.12U M=1 
X7 Y C1 net49 VSS LPNFET W=0.66U L=0.12U M=1 
X8 net49 A0 net55 VSS LPNFET W=0.66U L=0.12U M=1 
X9 net49 A1 net55 VSS LPNFET W=0.66U L=0.12U M=1 
.ENDS OAI222X1TS 

**** 
*.SUBCKT OAI222X2TS Y A0 A1 B0 B1 C0 C1 
.SUBCKT OAI222X2TS Y A0 A1 B0 B1 C0 C1 VSS VDD
X0 VDD B1 hnet18 VDD LPPFET W=0.84U L=0.12U M=1 
X1 hnet18 B0 Y VDD LPPFET W=0.84U L=0.12U M=1 
X10 VDD C1 hnet26 VDD LPPFET W=0.84U L=0.12U M=1 
X11 hnet26 C0 Y VDD LPPFET W=0.84U L=0.12U M=1 
X12 Y C0 net49 VSS LPNFET W=1.46U L=0.12U M=1 
X13 Y C1 net49 VSS LPNFET W=1.46U L=0.12U M=1 
X14 net49 A0 net55 VSS LPNFET W=1.46U L=0.12U M=1 
X15 net49 A1 net55 VSS LPNFET W=1.46U L=0.12U M=1 
X16 net55 B0 VSS VSS LPNFET W=1.32U L=0.12U M=1 
X17 net55 B1 VSS VSS LPNFET W=1.32U L=0.12U M=1 
X2 VDD B1 hnet14 VDD LPPFET W=0.84U L=0.12U M=1 
X3 hnet14 B0 Y VDD LPPFET W=0.84U L=0.12U M=1 
X4 VDD A1 hnet24 VDD LPPFET W=0.84U L=0.12U M=1 
X5 hnet24 A0 Y VDD LPPFET W=0.84U L=0.12U M=1 
X6 VDD A1 hnet20 VDD LPPFET W=0.84U L=0.12U M=1 
X7 hnet20 A0 Y VDD LPPFET W=0.84U L=0.12U M=1 
X8 VDD C1 hnet30 VDD LPPFET W=0.84U L=0.12U M=1 
X9 hnet30 C0 Y VDD LPPFET W=0.84U L=0.12U M=1 
.ENDS OAI222X2TS 

**** 
*.SUBCKT OAI222X4TS Y A0 A1 B0 B1 C0 C1 
.SUBCKT OAI222X4TS Y A0 A1 B0 B1 C0 C1 VSS VDD
X0 VDD net34 net30 VDD LPPFET W=1.02U L=0.12U M=1 
X1 net30 net34 VSS VSS LPNFET W=0.68U L=0.12U M=1 
X10 net34 C0 net54 VSS LPNFET W=0.46U L=0.12U M=1 
X11 net34 C1 net54 VSS LPNFET W=0.46U L=0.12U M=1 
X12 net54 A0 net60 VSS LPNFET W=0.46U L=0.12U M=1 
X13 net54 A1 net60 VSS LPNFET W=0.46U L=0.12U M=1 
X14 net60 B0 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X15 net60 B1 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X2 VDD net30 Y VDD LPPFET W=2.56U L=0.12U M=1 
X3 Y net30 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X4 VDD B1 hnet24 VDD LPPFET W=0.54U L=0.12U M=1 
X5 hnet24 B0 net34 VDD LPPFET W=0.54U L=0.12U M=1 
X6 VDD A1 hnet28 VDD LPPFET W=0.54U L=0.12U M=1 
X7 hnet28 A0 net34 VDD LPPFET W=0.54U L=0.12U M=1 
X8 VDD C1 hnet32 VDD LPPFET W=0.54U L=0.12U M=1 
X9 hnet32 C0 net34 VDD LPPFET W=0.54U L=0.12U M=1 
.ENDS OAI222X4TS 

**** 
*.SUBCKT OAI222XLTS Y A0 A1 B0 B1 C0 C1 
.SUBCKT OAI222XLTS Y A0 A1 B0 B1 C0 C1 VSS VDD
X0 VDD B1 hnet17 VDD LPPFET W=0.44U L=0.12U M=1 
X1 hnet17 B0 Y VDD LPPFET W=0.44U L=0.12U M=1 
X10 net55 B0 VSS VSS LPNFET W=0.48U L=0.12U M=1 
X11 net55 B1 VSS VSS LPNFET W=0.48U L=0.12U M=1 
X2 VDD A1 hnet22 VDD LPPFET W=0.44U L=0.12U M=1 
X3 hnet22 A0 Y VDD LPPFET W=0.44U L=0.12U M=1 
X4 VDD C1 hnet27 VDD LPPFET W=0.44U L=0.12U M=1 
X5 hnet27 C0 Y VDD LPPFET W=0.44U L=0.12U M=1 
X6 Y C0 net49 VSS LPNFET W=0.48U L=0.12U M=1 
X7 Y C1 net49 VSS LPNFET W=0.48U L=0.12U M=1 
X8 net49 A0 net55 VSS LPNFET W=0.48U L=0.12U M=1 
X9 net49 A1 net55 VSS LPNFET W=0.48U L=0.12U M=1 
.ENDS OAI222XLTS 

**** 
*.SUBCKT OAI22X1TS Y A0 A1 B0 B1 
.SUBCKT OAI22X1TS Y A0 A1 B0 B1 VSS VDD
X0 VDD B1 hnet14 VDD LPPFET W=0.84U L=0.12U M=1 
X1 hnet14 B0 Y VDD LPPFET W=0.84U L=0.12U M=1 
X2 VDD A1 hnet19 VDD LPPFET W=0.84U L=0.12U M=1 
X3 hnet19 A0 Y VDD LPPFET W=0.84U L=0.12U M=1 
X4 Y A0 net38 VSS LPNFET W=0.6U L=0.12U M=1 
X5 Y A1 net38 VSS LPNFET W=0.6U L=0.12U M=1 
X6 net38 B0 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X7 net38 B1 VSS VSS LPNFET W=0.6U L=0.12U M=1 
.ENDS OAI22X1TS 

**** 
*.SUBCKT OAI22X2TS Y A0 A1 B0 B1 
.SUBCKT OAI22X2TS Y A0 A1 B0 B1 VSS VDD
X0 VDD B1 hnet15 VDD LPPFET W=0.84U L=0.12U M=1 
X1 hnet15 B0 Y VDD LPPFET W=0.84U L=0.12U M=1 
X10 net38 B0 VSS VSS LPNFET W=1.22U L=0.12U M=1 
X11 net38 B1 VSS VSS LPNFET W=1.22U L=0.12U M=1 
X2 VDD B1 hnet11 VDD LPPFET W=0.84U L=0.12U M=1 
X3 hnet11 B0 Y VDD LPPFET W=0.84U L=0.12U M=1 
X4 VDD A1 hnet21 VDD LPPFET W=0.84U L=0.12U M=1 
X5 hnet21 A0 Y VDD LPPFET W=0.84U L=0.12U M=1 
X6 VDD A1 hnet17 VDD LPPFET W=0.84U L=0.12U M=1 
X7 hnet17 A0 Y VDD LPPFET W=0.84U L=0.12U M=1 
X8 Y A0 net38 VSS LPNFET W=1.22U L=0.12U M=1 
X9 Y A1 net38 VSS LPNFET W=1.22U L=0.12U M=1 
.ENDS OAI22X2TS 

**** 
*.SUBCKT OAI22X4TS Y A0 A1 B0 B1 
.SUBCKT OAI22X4TS Y A0 A1 B0 B1 VSS VDD
X0 VDD B1 hnet15 VDD LPPFET W=1.12U L=0.12U M=1 
X1 hnet15 B0 Y VDD LPPFET W=1.12U L=0.12U M=1 
X10 VDD A1 hnet17 VDD LPPFET W=1.12U L=0.12U M=1 
X11 hnet17 A0 Y VDD LPPFET W=1.12U L=0.12U M=1 
X12 Y A0 net38 VSS LPNFET W=2.44U L=0.12U M=1 
X13 Y A1 net38 VSS LPNFET W=2.44U L=0.12U M=1 
X14 net38 B0 VSS VSS LPNFET W=2.44U L=0.12U M=1 
X15 net38 B1 VSS VSS LPNFET W=2.44U L=0.12U M=1 
X2 VDD B1 hnet11 VDD LPPFET W=1.12U L=0.12U M=1 
X3 hnet11 B0 Y VDD LPPFET W=1.12U L=0.12U M=1 
X4 VDD B1 hnet10 VDD LPPFET W=1.12U L=0.12U M=1 
X5 hnet10 B0 Y VDD LPPFET W=1.12U L=0.12U M=1 
X6 VDD A1 hnet22 VDD LPPFET W=1.12U L=0.12U M=1 
X7 hnet22 A0 Y VDD LPPFET W=1.12U L=0.12U M=1 
X8 VDD A1 hnet18 VDD LPPFET W=1.12U L=0.12U M=1 
X9 hnet18 A0 Y VDD LPPFET W=1.12U L=0.12U M=1 
.ENDS OAI22X4TS 

**** 
*.SUBCKT OAI22XLTS Y A0 A1 B0 B1 
.SUBCKT OAI22XLTS Y A0 A1 B0 B1 VSS VDD
X0 VDD B1 hnet14 VDD LPPFET W=0.44U L=0.12U M=1 
X1 hnet14 B0 Y VDD LPPFET W=0.44U L=0.12U M=1 
X2 VDD A1 hnet19 VDD LPPFET W=0.44U L=0.12U M=1 
X3 hnet19 A0 Y VDD LPPFET W=0.44U L=0.12U M=1 
X4 Y A0 net38 VSS LPNFET W=0.4U L=0.12U M=1 
X5 Y A1 net38 VSS LPNFET W=0.4U L=0.12U M=1 
X6 net38 B0 VSS VSS LPNFET W=0.4U L=0.12U M=1 
X7 net38 B1 VSS VSS LPNFET W=0.4U L=0.12U M=1 
.ENDS OAI22XLTS 

**** 
*.SUBCKT OAI2BB1X1TS Y A0N A1N B0 
.SUBCKT OAI2BB1X1TS Y A0N A1N B0 VSS VDD
X0 hnet13 A0N VSS VSS LPNFET W=0.28U L=0.12U M=1 
X1 net11 A1N hnet13 VSS LPNFET W=0.28U L=0.12U M=1 
X2 VDD A0N net11 VDD LPPFET W=0.3U L=0.12U M=1 
X3 VDD A1N net11 VDD LPPFET W=0.3U L=0.12U M=1 
X4 hnet19 B0 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X5 Y net11 hnet19 VSS LPNFET W=0.6U L=0.12U M=1 
X6 VDD B0 Y VDD LPPFET W=0.64U L=0.12U M=1 
X7 VDD net11 Y VDD LPPFET W=0.64U L=0.12U M=1 
.ENDS OAI2BB1X1TS 

**** 
*.SUBCKT OAI2BB1X2TS Y A0N A1N B0 
.SUBCKT OAI2BB1X2TS Y A0N A1N B0 VSS VDD
X0 hnet13 A0N VSS VSS LPNFET W=0.54U L=0.12U M=1 
X1 net11 A1N hnet13 VSS LPNFET W=0.54U L=0.12U M=1 
X2 VDD A0N net11 VDD LPPFET W=0.56U L=0.12U M=1 
X3 VDD A1N net11 VDD LPPFET W=0.56U L=0.12U M=1 
X4 hnet18 B0 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X5 Y net11 hnet18 VSS LPNFET W=0.6U L=0.12U M=1 
X6 hnet14 B0 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X7 Y net11 hnet14 VSS LPNFET W=0.6U L=0.12U M=1 
X8 VDD B0 Y VDD LPPFET W=1.26U L=0.12U M=1 
X9 VDD net11 Y VDD LPPFET W=1.26U L=0.12U M=1 
.ENDS OAI2BB1X2TS 

**** 
*.SUBCKT OAI2BB1X4TS Y A0N A1N B0 
.SUBCKT OAI2BB1X4TS Y A0N A1N B0 VSS VDD
X0 hnet8 B0 VSS VSS LPNFET W=0.82U L=0.12U M=1 
X1 Y net14 hnet8 VSS LPNFET W=0.82U L=0.12U M=1 
X10 VDD A0N net14 VDD LPPFET W=1.06U L=0.12U M=1 
X11 VDD A1N net14 VDD LPPFET W=1.06U L=0.12U M=1 
X2 hnet9 B0 VSS VSS LPNFET W=0.82U L=0.12U M=1 
X3 Y net14 hnet9 VSS LPNFET W=0.82U L=0.12U M=1 
X4 hnet12 B0 VSS VSS LPNFET W=0.82U L=0.12U M=1 
X5 Y net14 hnet12 VSS LPNFET W=0.82U L=0.12U M=1 
X6 VDD B0 Y VDD LPPFET W=2.56U L=0.12U M=1 
X7 VDD net14 Y VDD LPPFET W=2.56U L=0.12U M=1 
X8 hnet19 A0N VSS VSS LPNFET W=0.84U L=0.12U M=1 
X9 net14 A1N hnet19 VSS LPNFET W=0.84U L=0.12U M=1 
.ENDS OAI2BB1X4TS 

**** 
*.SUBCKT OAI2BB1XLTS Y A0N A1N B0 
.SUBCKT OAI2BB1XLTS Y A0N A1N B0 VSS VDD
X0 hnet13 A0N VSS VSS LPNFET W=0.26U L=0.12U M=1 
X1 net11 A1N hnet13 VSS LPNFET W=0.26U L=0.12U M=1 
X2 VDD A0N net11 VDD LPPFET W=0.28U L=0.12U M=1 
X3 VDD A1N net11 VDD LPPFET W=0.28U L=0.12U M=1 
X4 hnet19 B0 VSS VSS LPNFET W=0.4U L=0.12U M=1 
X5 Y net11 hnet19 VSS LPNFET W=0.4U L=0.12U M=1 
X6 VDD B0 Y VDD LPPFET W=0.42U L=0.12U M=1 
X7 VDD net11 Y VDD LPPFET W=0.42U L=0.12U M=1 
.ENDS OAI2BB1XLTS 

**** 
*.SUBCKT OAI2BB2X1TS Y A0N A1N B0 B1 
.SUBCKT OAI2BB2X1TS Y A0N A1N B0 B1 VSS VDD
X0 VDD B1 hnet15 VDD LPPFET W=0.84U L=0.12U M=1 
X1 hnet15 B0 Y VDD LPPFET W=0.84U L=0.12U M=1 
X2 hnet19 A0N VSS VSS LPNFET W=0.28U L=0.12U M=1 
X3 nmin1 A1N hnet19 VSS LPNFET W=0.28U L=0.12U M=1 
X4 VDD A0N nmin1 VDD LPPFET W=0.3U L=0.12U M=1 
X5 VDD A1N nmin1 VDD LPPFET W=0.3U L=0.12U M=1 
X6 Y nmin1 VDD VDD LPPFET W=0.64U L=0.12U M=1 
X7 net33 B0 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X8 Y nmin1 net33 VSS LPNFET W=0.6U L=0.12U M=1 
X9 net33 B1 VSS VSS LPNFET W=0.6U L=0.12U M=1 
.ENDS OAI2BB2X1TS 

**** 
*.SUBCKT OAI2BB2X2TS Y A0N A1N B0 B1 
.SUBCKT OAI2BB2X2TS Y A0N A1N B0 B1 VSS VDD
X0 VDD B1 hnet16 VDD LPPFET W=0.84U L=0.12U M=1 
X1 hnet16 B0 Y VDD LPPFET W=0.84U L=0.12U M=1 
X10 Y nmin1 net33 VSS LPNFET W=1.22U L=0.12U M=1 
X11 net33 B1 VSS VSS LPNFET W=1.22U L=0.12U M=1 
X2 VDD B1 hnet13 VDD LPPFET W=0.84U L=0.12U M=1 
X3 hnet13 B0 Y VDD LPPFET W=0.84U L=0.12U M=1 
X4 hnet20 A0N VSS VSS LPNFET W=0.56U L=0.12U M=1 
X5 nmin1 A1N hnet20 VSS LPNFET W=0.56U L=0.12U M=1 
X6 VDD A0N nmin1 VDD LPPFET W=0.58U L=0.12U M=1 
X7 VDD A1N nmin1 VDD LPPFET W=0.58U L=0.12U M=1 
X8 Y nmin1 VDD VDD LPPFET W=1.28U L=0.12U M=1 
X9 net33 B0 VSS VSS LPNFET W=1.22U L=0.12U M=1 
.ENDS OAI2BB2X2TS 

**** 
*.SUBCKT OAI2BB2X4TS Y A0N A1N B0 B1 
.SUBCKT OAI2BB2X4TS Y A0N A1N B0 B1 VSS VDD
X0 VDD B1 hnet16 VDD LPPFET W=1.12U L=0.12U M=1 
X1 hnet16 B0 Y VDD LPPFET W=1.12U L=0.12U M=1 
X10 Y nmin1 VDD VDD LPPFET W=2.56U L=0.12U M=1 
X11 net33 B0 VSS VSS LPNFET W=2.44U L=0.12U M=1 
X12 Y nmin1 net33 VSS LPNFET W=2.42U L=0.12U M=1 
X13 net33 B1 VSS VSS LPNFET W=2.44U L=0.12U M=1 
X2 VDD B1 hnet13 VDD LPPFET W=1.12U L=0.12U M=1 
X3 hnet13 B0 Y VDD LPPFET W=1.12U L=0.12U M=1 
X4 VDD B1 hnet12 VDD LPPFET W=1.12U L=0.12U M=1 
X5 hnet12 B0 Y VDD LPPFET W=1.12U L=0.12U M=1 
X6 hnet21 A0N VSS VSS LPNFET W=0.92U L=0.12U M=1 
X7 nmin1 A1N hnet21 VSS LPNFET W=0.92U L=0.12U M=1 
X8 VDD A0N nmin1 VDD LPPFET W=1.18U L=0.12U M=1 
X9 VDD A1N nmin1 VDD LPPFET W=1.18U L=0.12U M=1 
.ENDS OAI2BB2X4TS 

**** 
*.SUBCKT OAI2BB2XLTS Y A0N A1N B0 B1 
.SUBCKT OAI2BB2XLTS Y A0N A1N B0 B1 VSS VDD
X0 VDD B1 hnet15 VDD LPPFET W=0.44U L=0.12U M=1 
X1 hnet15 B0 Y VDD LPPFET W=0.44U L=0.12U M=1 
X2 hnet19 A0N VSS VSS LPNFET W=0.26U L=0.12U M=1 
X3 nmin1 A1N hnet19 VSS LPNFET W=0.26U L=0.12U M=1 
X4 VDD A0N nmin1 VDD LPPFET W=0.28U L=0.12U M=1 
X5 VDD A1N nmin1 VDD LPPFET W=0.28U L=0.12U M=1 
X6 Y nmin1 VDD VDD LPPFET W=0.42U L=0.12U M=1 
X7 net33 B0 VSS VSS LPNFET W=0.4U L=0.12U M=1 
X8 Y nmin1 net33 VSS LPNFET W=0.4U L=0.12U M=1 
X9 net33 B1 VSS VSS LPNFET W=0.4U L=0.12U M=1 
.ENDS OAI2BB2XLTS 

**** 
*.SUBCKT OAI31X1TS Y A0 A1 A2 B0 
.SUBCKT OAI31X1TS Y A0 A1 A2 B0 VSS VDD
X0 VDD A2 hnet11 VDD LPPFET W=1.02U L=0.12U M=1 
X1 hnet11 A1 hnet16 VDD LPPFET W=1.02U L=0.12U M=1 
X2 hnet16 A0 Y VDD LPPFET W=1.02U L=0.12U M=1 
X3 net24 A0 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X4 Y B0 net24 VSS LPNFET W=0.6U L=0.12U M=1 
X5 net24 A2 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X6 net24 A1 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X7 Y B0 VDD VDD LPPFET W=0.64U L=0.12U M=1 
.ENDS OAI31X1TS 

**** 
*.SUBCKT OAI31X2TS Y A0 A1 A2 B0 
.SUBCKT OAI31X2TS Y A0 A1 A2 B0 VSS VDD
X0 VDD A2 hnet12 VDD LPPFET W=1.04U L=0.12U M=1 
X1 hnet12 A1 hnet11 VDD LPPFET W=1.04U L=0.12U M=1 
X10 Y B0 VDD VDD LPPFET W=1.28U L=0.12U M=1 
X2 hnet11 A0 Y VDD LPPFET W=1.04U L=0.12U M=1 
X3 VDD A2 hnet14 VDD LPPFET W=1.04U L=0.12U M=1 
X4 hnet14 A1 hnet15 VDD LPPFET W=1.04U L=0.12U M=1 
X5 hnet15 A0 Y VDD LPPFET W=1.04U L=0.12U M=1 
X6 net24 A0 VSS VSS LPNFET W=1.22U L=0.12U M=1 
X7 Y B0 net24 VSS LPNFET W=1.22U L=0.12U M=1 
X8 net24 A2 VSS VSS LPNFET W=1.22U L=0.12U M=1 
X9 net24 A1 VSS VSS LPNFET W=1.22U L=0.12U M=1 
.ENDS OAI31X2TS 

**** 
*.SUBCKT OAI31X4TS Y A0 A1 A2 B0 
.SUBCKT OAI31X4TS Y A0 A1 A2 B0 VSS VDD
X0 VDD net23 net19 VDD LPPFET W=1.02U L=0.12U M=1 
X1 net19 net23 VSS VSS LPNFET W=0.74U L=0.12U M=1 
X10 net29 A1 VSS VSS LPNFET W=0.38U L=0.12U M=1 
X11 net23 B0 VDD VDD LPPFET W=0.4U L=0.12U M=1 
X2 VDD net19 Y VDD LPPFET W=2.56U L=0.12U M=1 
X3 Y net19 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X4 VDD A2 hnet17 VDD LPPFET W=0.66U L=0.12U M=1 
X5 hnet17 A1 hnet22 VDD LPPFET W=0.66U L=0.12U M=1 
X6 hnet22 A0 net23 VDD LPPFET W=0.66U L=0.12U M=1 
X7 net29 A0 VSS VSS LPNFET W=0.38U L=0.12U M=1 
X8 net23 B0 net29 VSS LPNFET W=0.38U L=0.12U M=1 
X9 net29 A2 VSS VSS LPNFET W=0.38U L=0.12U M=1 
.ENDS OAI31X4TS 

**** 
*.SUBCKT OAI31XLTS Y A0 A1 A2 B0 
.SUBCKT OAI31XLTS Y A0 A1 A2 B0 VSS VDD
X0 VDD A2 hnet11 VDD LPPFET W=0.54U L=0.12U M=1 
X1 hnet11 A1 hnet16 VDD LPPFET W=0.54U L=0.12U M=1 
X2 hnet16 A0 Y VDD LPPFET W=0.54U L=0.12U M=1 
X3 net24 A0 VSS VSS LPNFET W=0.4U L=0.12U M=1 
X4 Y B0 net24 VSS LPNFET W=0.4U L=0.12U M=1 
X5 net24 A2 VSS VSS LPNFET W=0.4U L=0.12U M=1 
X6 net24 A1 VSS VSS LPNFET W=0.4U L=0.12U M=1 
X7 Y B0 VDD VDD LPPFET W=0.42U L=0.12U M=1 
.ENDS OAI31XLTS 

**** 
*.SUBCKT OAI32X1TS Y A0 A1 A2 B0 B1 
.SUBCKT OAI32X1TS Y A0 A1 A2 B0 B1 VSS VDD
X0 VDD A2 hnet11 VDD LPPFET W=1.02U L=0.12U M=1 
X1 hnet11 A1 hnet17 VDD LPPFET W=1.02U L=0.12U M=1 
X2 hnet17 A0 Y VDD LPPFET W=1.02U L=0.12U M=1 
X3 VDD B1 hnet21 VDD LPPFET W=0.84U L=0.12U M=1 
X4 hnet21 B0 Y VDD LPPFET W=0.84U L=0.12U M=1 
X5 net46 A0 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X6 Y B0 net46 VSS LPNFET W=0.6U L=0.12U M=1 
X7 Y B1 net46 VSS LPNFET W=0.6U L=0.12U M=1 
X8 net46 A1 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X9 net46 A2 VSS VSS LPNFET W=0.6U L=0.12U M=1 
.ENDS OAI32X1TS 

**** 
*.SUBCKT OAI32X2TS Y A0 A1 A2 B0 B1 
.SUBCKT OAI32X2TS Y A0 A1 A2 B0 B1 VSS VDD
X0 VDD A2 hnet12 VDD LPPFET W=1.04U L=0.12U M=1 
X1 hnet12 A1 hnet11 VDD LPPFET W=1.04U L=0.12U M=1 
X10 net46 A0 VSS VSS LPNFET W=1.22U L=0.12U M=1 
X11 Y B0 net46 VSS LPNFET W=1.16U L=0.12U M=1 
X12 Y B1 net46 VSS LPNFET W=1.16U L=0.12U M=1 
X13 net46 A1 VSS VSS LPNFET W=1.22U L=0.12U M=1 
X14 net46 A2 VSS VSS LPNFET W=1.22U L=0.12U M=1 
X2 hnet11 A0 Y VDD LPPFET W=1.04U L=0.12U M=1 
X3 VDD A2 hnet14 VDD LPPFET W=1.04U L=0.12U M=1 
X4 hnet14 A1 hnet15 VDD LPPFET W=1.04U L=0.12U M=1 
X5 hnet15 A0 Y VDD LPPFET W=1.04U L=0.12U M=1 
X6 VDD B1 hnet24 VDD LPPFET W=0.84U L=0.12U M=1 
X7 hnet24 B0 Y VDD LPPFET W=0.84U L=0.12U M=1 
X8 VDD B1 hnet21 VDD LPPFET W=0.84U L=0.12U M=1 
X9 hnet21 B0 Y VDD LPPFET W=0.84U L=0.12U M=1 
.ENDS OAI32X2TS 

**** 
*.SUBCKT OAI32X4TS Y A0 A1 A2 B0 B1 
.SUBCKT OAI32X4TS Y A0 A1 A2 B0 B1 VSS VDD
X0 VDD net26 net22 VDD LPPFET W=1.02U L=0.12U M=1 
X1 net22 net26 VSS VSS LPNFET W=0.74U L=0.12U M=1 
X10 net26 B0 net47 VSS LPNFET W=0.38U L=0.12U M=1 
X11 net26 B1 net47 VSS LPNFET W=0.38U L=0.12U M=1 
X12 net47 A1 VSS VSS LPNFET W=0.38U L=0.12U M=1 
X13 net47 A2 VSS VSS LPNFET W=0.38U L=0.12U M=1 
X2 VDD net22 Y VDD LPPFET W=2.56U L=0.12U M=1 
X3 Y net22 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X4 VDD A2 hnet19 VDD LPPFET W=0.66U L=0.12U M=1 
X5 hnet19 A1 hnet24 VDD LPPFET W=0.66U L=0.12U M=1 
X6 hnet24 A0 net26 VDD LPPFET W=0.66U L=0.12U M=1 
X7 VDD B1 hnet28 VDD LPPFET W=0.54U L=0.12U M=1 
X8 hnet28 B0 net26 VDD LPPFET W=0.54U L=0.12U M=1 
X9 net47 A0 VSS VSS LPNFET W=0.38U L=0.12U M=1 
.ENDS OAI32X4TS 

**** 
*.SUBCKT OAI32XLTS Y A0 A1 A2 B0 B1 
.SUBCKT OAI32XLTS Y A0 A1 A2 B0 B1 VSS VDD
X0 VDD A2 hnet11 VDD LPPFET W=0.54U L=0.12U M=1 
X1 hnet11 A1 hnet17 VDD LPPFET W=0.54U L=0.12U M=1 
X2 hnet17 A0 Y VDD LPPFET W=0.54U L=0.12U M=1 
X3 VDD B1 hnet21 VDD LPPFET W=0.44U L=0.12U M=1 
X4 hnet21 B0 Y VDD LPPFET W=0.44U L=0.12U M=1 
X5 net46 A0 VSS VSS LPNFET W=0.4U L=0.12U M=1 
X6 Y B0 net46 VSS LPNFET W=0.4U L=0.12U M=1 
X7 Y B1 net46 VSS LPNFET W=0.4U L=0.12U M=1 
X8 net46 A1 VSS VSS LPNFET W=0.4U L=0.12U M=1 
X9 net46 A2 VSS VSS LPNFET W=0.4U L=0.12U M=1 
.ENDS OAI32XLTS 

**** 
*.SUBCKT OAI33X1TS Y A0 A1 A2 B0 B1 B2 
.SUBCKT OAI33X1TS Y A0 A1 A2 B0 B1 B2 VSS VDD
X0 VDD A2 hnet12 VDD LPPFET W=1.02U L=0.12U M=1 
X1 hnet12 A1 hnet18 VDD LPPFET W=1.02U L=0.12U M=1 
X10 net57 B1 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X11 net57 B2 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X2 hnet18 A0 Y VDD LPPFET W=1.02U L=0.12U M=1 
X3 VDD B2 hnet19 VDD LPPFET W=1.02U L=0.12U M=1 
X4 hnet19 B1 hnet25 VDD LPPFET W=1.02U L=0.12U M=1 
X5 hnet25 B0 Y VDD LPPFET W=1.02U L=0.12U M=1 
X6 net57 B0 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X7 Y A0 net57 VSS LPNFET W=0.6U L=0.12U M=1 
X8 Y A1 net57 VSS LPNFET W=0.6U L=0.12U M=1 
X9 Y A2 net57 VSS LPNFET W=0.6U L=0.12U M=1 
.ENDS OAI33X1TS 

**** 
*.SUBCKT OAI33X2TS Y A0 A1 A2 B0 B1 B2 
.SUBCKT OAI33X2TS Y A0 A1 A2 B0 B1 B2 VSS VDD
X0 VDD A2 hnet13 VDD LPPFET W=1.04U L=0.12U M=1 
X1 hnet13 A1 hnet12 VDD LPPFET W=1.04U L=0.12U M=1 
X10 hnet24 B1 hnet25 VDD LPPFET W=1.04U L=0.12U M=1 
X11 hnet25 B0 Y VDD LPPFET W=1.04U L=0.12U M=1 
X12 net57 B0 VSS VSS LPNFET W=1.22U L=0.12U M=1 
X13 Y A0 net57 VSS LPNFET W=1.16U L=0.12U M=1 
X14 Y A1 net57 VSS LPNFET W=1.16U L=0.12U M=1 
X15 Y A2 net57 VSS LPNFET W=1.16U L=0.12U M=1 
X16 net57 B1 VSS VSS LPNFET W=1.22U L=0.12U M=1 
X17 net57 B2 VSS VSS LPNFET W=1.22U L=0.12U M=1 
X2 hnet12 A0 Y VDD LPPFET W=1.04U L=0.12U M=1 
X3 VDD A2 hnet15 VDD LPPFET W=1.04U L=0.12U M=1 
X4 hnet15 A1 hnet16 VDD LPPFET W=1.04U L=0.12U M=1 
X5 hnet16 A0 Y VDD LPPFET W=1.04U L=0.12U M=1 
X6 VDD B2 hnet22 VDD LPPFET W=1.04U L=0.12U M=1 
X7 hnet22 B1 hnet21 VDD LPPFET W=1.04U L=0.12U M=1 
X8 hnet21 B0 Y VDD LPPFET W=1.04U L=0.12U M=1 
X9 VDD B2 hnet24 VDD LPPFET W=1.04U L=0.12U M=1 
.ENDS OAI33X2TS 

**** 
*.SUBCKT OAI33X4TS Y A0 A1 A2 B0 B1 B2 
.SUBCKT OAI33X4TS Y A0 A1 A2 B0 B1 B2 VSS VDD
X0 VDD net41 net33 VDD LPPFET W=1.02U L=0.12U M=1 
X1 net33 net41 VSS VSS LPNFET W=0.74U L=0.12U M=1 
X10 net62 B0 VSS VSS LPNFET W=0.38U L=0.12U M=1 
X11 net41 A0 net62 VSS LPNFET W=0.38U L=0.12U M=1 
X12 net41 A1 net62 VSS LPNFET W=0.38U L=0.12U M=1 
X13 net41 A2 net62 VSS LPNFET W=0.38U L=0.12U M=1 
X14 net62 B1 VSS VSS LPNFET W=0.38U L=0.12U M=1 
X15 net62 B2 VSS VSS LPNFET W=0.38U L=0.12U M=1 
X2 VDD net33 Y VDD LPPFET W=2.48U L=0.12U M=1 
X3 Y net33 VSS VSS LPNFET W=1.78U L=0.12U M=1 
X4 VDD A2 hnet20 VDD LPPFET W=0.66U L=0.12U M=1 
X5 hnet20 A1 hnet25 VDD LPPFET W=0.66U L=0.12U M=1 
X6 hnet25 A0 net41 VDD LPPFET W=0.66U L=0.12U M=1 
X7 VDD B2 hnet26 VDD LPPFET W=0.66U L=0.12U M=1 
X8 hnet26 B1 hnet31 VDD LPPFET W=0.66U L=0.12U M=1 
X9 hnet31 B0 net41 VDD LPPFET W=0.66U L=0.12U M=1 
.ENDS OAI33X4TS 

**** 
*.SUBCKT OAI33XLTS Y A0 A1 A2 B0 B1 B2 
.SUBCKT OAI33XLTS Y A0 A1 A2 B0 B1 B2 VSS VDD
X0 VDD A2 hnet12 VDD LPPFET W=0.54U L=0.12U M=1 
X1 hnet12 A1 hnet18 VDD LPPFET W=0.54U L=0.12U M=1 
X10 net57 B1 VSS VSS LPNFET W=0.4U L=0.12U M=1 
X11 net57 B2 VSS VSS LPNFET W=0.4U L=0.12U M=1 
X2 hnet18 A0 Y VDD LPPFET W=0.54U L=0.12U M=1 
X3 VDD B2 hnet19 VDD LPPFET W=0.54U L=0.12U M=1 
X4 hnet19 B1 hnet25 VDD LPPFET W=0.54U L=0.12U M=1 
X5 hnet25 B0 Y VDD LPPFET W=0.54U L=0.12U M=1 
X6 net57 B0 VSS VSS LPNFET W=0.4U L=0.12U M=1 
X7 Y A0 net57 VSS LPNFET W=0.4U L=0.12U M=1 
X8 Y A1 net57 VSS LPNFET W=0.4U L=0.12U M=1 
X9 Y A2 net57 VSS LPNFET W=0.4U L=0.12U M=1 
.ENDS OAI33XLTS 

**** 
*.SUBCKT OR2X1TS Y A B 
.SUBCKT OR2X1TS Y A B VSS VDD
X0 VDD nmin Y VDD LPPFET W=0.64U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=0.46U L=0.12U M=1 
X2 nmin B VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 nmin A VSS VSS LPNFET W=0.2U L=0.12U M=1 
X4 VDD B hnet12 VDD LPPFET W=0.36U L=0.12U M=1 
X5 hnet12 A nmin VDD LPPFET W=0.36U L=0.12U M=1 
.ENDS OR2X1TS 

**** 
*.SUBCKT OR2X2TS Y A B 
.SUBCKT OR2X2TS Y A B VSS VDD
X0 VDD nmin Y VDD LPPFET W=1.28U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=0.92U L=0.12U M=1 
X2 nmin B VSS VSS LPNFET W=0.36U L=0.12U M=1 
X3 nmin A VSS VSS LPNFET W=0.36U L=0.12U M=1 
X4 VDD B hnet12 VDD LPPFET W=0.66U L=0.12U M=1 
X5 hnet12 A nmin VDD LPPFET W=0.66U L=0.12U M=1 
.ENDS OR2X2TS 

**** 
*.SUBCKT OR2X4TS Y A B 
.SUBCKT OR2X4TS Y A B VSS VDD
X0 VDD nmin Y VDD LPPFET W=2.46U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=1.84U L=0.12U M=1 
X2 nmin B VSS VSS LPNFET W=0.66U L=0.12U M=1 
X3 nmin A VSS VSS LPNFET W=0.66U L=0.12U M=1 
X4 VDD B hnet12 VDD LPPFET W=1.3U L=0.12U M=1 
X5 hnet12 A nmin VDD LPPFET W=1.3U L=0.12U M=1 
.ENDS OR2X4TS 

**** 
*.SUBCKT OR2X6TS Y A B 
.SUBCKT OR2X6TS Y A B VSS VDD
X0 VDD nmin Y VDD LPPFET W=3.84U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=2.76U L=0.12U M=1 
X2 nmin B VSS VSS LPNFET W=1.1U L=0.12U M=1 
X3 nmin A VSS VSS LPNFET W=1.1U L=0.12U M=1 
X4 VDD B hnet13 VDD LPPFET W=1U L=0.12U M=1 
X5 hnet13 A nmin VDD LPPFET W=1U L=0.12U M=1 
X6 VDD B hnet11 VDD LPPFET W=1U L=0.12U M=1 
X7 hnet11 A nmin VDD LPPFET W=1U L=0.12U M=1 
.ENDS OR2X6TS 

**** 
*.SUBCKT OR2X8TS Y A B 
.SUBCKT OR2X8TS Y A B VSS VDD
X0 VDD nmin Y VDD LPPFET W=4.68U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=3.42U L=0.12U M=1 
X2 nmin B VSS VSS LPNFET W=1.32U L=0.12U M=1 
X3 nmin A VSS VSS LPNFET W=1.32U L=0.12U M=1 
X4 VDD B hnet13 VDD LPPFET W=1.3U L=0.12U M=1 
X5 hnet13 A nmin VDD LPPFET W=1.3U L=0.12U M=1 
X6 VDD B hnet11 VDD LPPFET W=1.3U L=0.12U M=1 
X7 hnet11 A nmin VDD LPPFET W=1.3U L=0.12U M=1 
.ENDS OR2X8TS 

**** 
*.SUBCKT OR2XLTS A B Y 
.SUBCKT OR2XLTS A B Y VSS VDD
X0 VDD nmin Y VDD LPPFET W=0.42U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=0.24U L=0.12U M=1 
X2 nmin B VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 nmin A VSS VSS LPNFET W=0.2U L=0.12U M=1 
X4 VDD B hnet12 VDD LPPFET W=0.3U L=0.12U M=1 
X5 hnet12 A nmin VDD LPPFET W=0.3U L=0.12U M=1 
.ENDS OR2XLTS 

**** 
*.SUBCKT OR3X1TS Y A B C 
.SUBCKT OR3X1TS Y A B C VSS VDD
X0 VDD nmin Y VDD LPPFET W=0.64U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=0.46U L=0.12U M=1 
X2 nmin C VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 nmin B VSS VSS LPNFET W=0.2U L=0.12U M=1 
X4 nmin A VSS VSS LPNFET W=0.2U L=0.12U M=1 
X5 VDD C hnet17 VDD LPPFET W=0.44U L=0.12U M=1 
X6 hnet17 B hnet16 VDD LPPFET W=0.44U L=0.12U M=1 
X7 hnet16 A nmin VDD LPPFET W=0.44U L=0.12U M=1 
.ENDS OR3X1TS 

**** 
*.SUBCKT OR3X2TS Y A B C 
.SUBCKT OR3X2TS Y A B C VSS VDD
X0 VDD nmin Y VDD LPPFET W=1.28U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=0.92U L=0.12U M=1 
X2 nmin C VSS VSS LPNFET W=0.36U L=0.12U M=1 
X3 nmin B VSS VSS LPNFET W=0.36U L=0.12U M=1 
X4 nmin A VSS VSS LPNFET W=0.36U L=0.12U M=1 
X5 VDD C hnet17 VDD LPPFET W=0.8U L=0.12U M=1 
X6 hnet17 B hnet16 VDD LPPFET W=0.8U L=0.12U M=1 
X7 hnet16 A nmin VDD LPPFET W=0.8U L=0.12U M=1 
.ENDS OR3X2TS 

**** 
*.SUBCKT OR3X4TS Y A B C 
.SUBCKT OR3X4TS Y A B C VSS VDD
X0 VDD nmin Y VDD LPPFET W=2.56U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=1.84U L=0.12U M=1 
X10 hnet12 A nmin VDD LPPFET W=0.84U L=0.12U M=1 
X2 nmin C VSS VSS LPNFET W=0.74U L=0.12U M=1 
X3 nmin B VSS VSS LPNFET W=0.74U L=0.12U M=1 
X4 nmin A VSS VSS LPNFET W=0.74U L=0.12U M=1 
X5 VDD C hnet19 VDD LPPFET W=0.84U L=0.12U M=1 
X6 hnet19 B hnet15 VDD LPPFET W=0.84U L=0.12U M=1 
X7 hnet15 A nmin VDD LPPFET W=0.84U L=0.12U M=1 
X8 VDD C hnet14 VDD LPPFET W=0.84U L=0.12U M=1 
X9 hnet14 B hnet12 VDD LPPFET W=0.84U L=0.12U M=1 
.ENDS OR3X4TS 

**** 
*.SUBCKT OR3X6TS Y A B C 
.SUBCKT OR3X6TS Y A B C VSS VDD
X0 VDD nmin Y VDD LPPFET W=3.5U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=2.76U L=0.12U M=1 
X10 hnet12 A nmin VDD LPPFET W=1.24U L=0.12U M=1 
X2 nmin C VSS VSS LPNFET W=0.92U L=0.12U M=1 
X3 nmin B VSS VSS LPNFET W=0.92U L=0.12U M=1 
X4 nmin A VSS VSS LPNFET W=0.92U L=0.12U M=1 
X5 VDD C hnet19 VDD LPPFET W=1.24U L=0.12U M=1 
X6 hnet19 B hnet15 VDD LPPFET W=1.24U L=0.12U M=1 
X7 hnet15 A nmin VDD LPPFET W=1.24U L=0.12U M=1 
X8 VDD C hnet14 VDD LPPFET W=1.24U L=0.12U M=1 
X9 hnet14 B hnet12 VDD LPPFET W=1.24U L=0.12U M=1 
.ENDS OR3X6TS 

**** 
*.SUBCKT OR3X8TS Y A B C 
.SUBCKT OR3X8TS Y A B C VSS VDD
X0 VDD nmin Y VDD LPPFET W=5.12U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=3.68U L=0.12U M=1 
X10 hnet15 A nmin VDD LPPFET W=1.06U L=0.12U M=1 
X11 VDD C hnet12 VDD LPPFET W=1.06U L=0.12U M=1 
X12 hnet12 B hnet20 VDD LPPFET W=1.06U L=0.12U M=1 
X13 hnet20 A nmin VDD LPPFET W=1.06U L=0.12U M=1 
X2 nmin C VSS VSS LPNFET W=1.48U L=0.12U M=1 
X3 nmin B VSS VSS LPNFET W=1.48U L=0.12U M=1 
X4 nmin A VSS VSS LPNFET W=1.48U L=0.12U M=1 
X5 VDD C hnet21 VDD LPPFET W=1.06U L=0.12U M=1 
X6 hnet21 B hnet16 VDD LPPFET W=1.06U L=0.12U M=1 
X7 hnet16 A nmin VDD LPPFET W=1.06U L=0.12U M=1 
X8 VDD C hnet14 VDD LPPFET W=1.06U L=0.12U M=1 
X9 hnet14 B hnet15 VDD LPPFET W=1.06U L=0.12U M=1 
.ENDS OR3X8TS 

**** 
*.SUBCKT OR3XLTS Y A B C 
.SUBCKT OR3XLTS Y A B C VSS VDD
X0 VDD nmin Y VDD LPPFET W=0.42U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=0.24U L=0.12U M=1 
X2 nmin C VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 nmin B VSS VSS LPNFET W=0.2U L=0.12U M=1 
X4 nmin A VSS VSS LPNFET W=0.2U L=0.12U M=1 
X5 VDD C hnet17 VDD LPPFET W=0.36U L=0.12U M=1 
X6 hnet17 B hnet16 VDD LPPFET W=0.36U L=0.12U M=1 
X7 hnet16 A nmin VDD LPPFET W=0.36U L=0.12U M=1 
.ENDS OR3XLTS 

**** 
*.SUBCKT OR4X1TS Y A B C D 
.SUBCKT OR4X1TS Y A B C D VSS VDD
X0 VDD nmin Y VDD LPPFET W=0.64U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=0.46U L=0.12U M=1 
X2 nmin D VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 nmin C VSS VSS LPNFET W=0.2U L=0.12U M=1 
X4 nmin B VSS VSS LPNFET W=0.2U L=0.12U M=1 
X5 nmin A VSS VSS LPNFET W=0.2U L=0.12U M=1 
X6 VDD D hnet15 VDD LPPFET W=0.52U L=0.12U M=1 
X7 hnet15 C hnet18 VDD LPPFET W=0.52U L=0.12U M=1 
X8 hnet18 B hnet14 VDD LPPFET W=0.52U L=0.12U M=1 
X9 hnet14 A nmin VDD LPPFET W=0.52U L=0.12U M=1 
.ENDS OR4X1TS 

**** 
*.SUBCKT OR4X2TS Y A B C D 
.SUBCKT OR4X2TS Y A B C D VSS VDD
X0 VDD nmin Y VDD LPPFET W=1.28U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=0.92U L=0.12U M=1 
X2 nmin D VSS VSS LPNFET W=0.36U L=0.12U M=1 
X3 nmin C VSS VSS LPNFET W=0.36U L=0.12U M=1 
X4 nmin B VSS VSS LPNFET W=0.36U L=0.12U M=1 
X5 nmin A VSS VSS LPNFET W=0.36U L=0.12U M=1 
X6 VDD D hnet15 VDD LPPFET W=0.94U L=0.12U M=1 
X7 hnet15 C hnet18 VDD LPPFET W=0.94U L=0.12U M=1 
X8 hnet18 B hnet14 VDD LPPFET W=0.94U L=0.12U M=1 
X9 hnet14 A nmin VDD LPPFET W=0.94U L=0.12U M=1 
.ENDS OR4X2TS 

**** 
*.SUBCKT OR4X4TS Y A B C D 
.SUBCKT OR4X4TS Y A B C D VSS VDD
X0 VDD nmin Y VDD LPPFET W=2.56U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=1.84U L=0.12U M=1 
X10 VDD D hnet14 VDD LPPFET W=0.96U L=0.12U M=1 
X11 hnet14 C hnet13 VDD LPPFET W=0.96U L=0.12U M=1 
X12 hnet13 B hnet22 VDD LPPFET W=0.96U L=0.12U M=1 
X13 hnet22 A nmin VDD LPPFET W=0.96U L=0.12U M=1 
X2 nmin D VSS VSS LPNFET W=0.74U L=0.12U M=1 
X3 nmin C VSS VSS LPNFET W=0.74U L=0.12U M=1 
X4 nmin B VSS VSS LPNFET W=0.74U L=0.12U M=1 
X5 nmin A VSS VSS LPNFET W=0.74U L=0.12U M=1 
X6 VDD D hnet18 VDD LPPFET W=0.96U L=0.12U M=1 
X7 hnet18 C hnet17 VDD LPPFET W=0.96U L=0.12U M=1 
X8 hnet17 B hnet16 VDD LPPFET W=0.96U L=0.12U M=1 
X9 hnet16 A nmin VDD LPPFET W=0.96U L=0.12U M=1 
.ENDS OR4X4TS 

**** 
*.SUBCKT OR4X6TS Y A B C D 
.SUBCKT OR4X6TS Y A B C D VSS VDD
X0 VDD nmin Y VDD LPPFET W=3.64U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=2.76U L=0.12U M=1 
X10 VDD D hnet14 VDD LPPFET W=1.3U L=0.12U M=1 
X11 hnet14 C hnet13 VDD LPPFET W=1.3U L=0.12U M=1 
X12 hnet13 B hnet22 VDD LPPFET W=1.3U L=0.12U M=1 
X13 hnet22 A nmin VDD LPPFET W=1.3U L=0.12U M=1 
X2 nmin D VSS VSS LPNFET W=1.08U L=0.12U M=1 
X3 nmin C VSS VSS LPNFET W=1.08U L=0.12U M=1 
X4 nmin B VSS VSS LPNFET W=1.08U L=0.12U M=1 
X5 nmin A VSS VSS LPNFET W=1.08U L=0.12U M=1 
X6 VDD D hnet18 VDD LPPFET W=1.3U L=0.12U M=1 
X7 hnet18 C hnet17 VDD LPPFET W=1.3U L=0.12U M=1 
X8 hnet17 B hnet16 VDD LPPFET W=1.3U L=0.12U M=1 
X9 hnet16 A nmin VDD LPPFET W=1.3U L=0.12U M=1 
.ENDS OR4X6TS 

**** 
*.SUBCKT OR4X8TS Y A B C D 
.SUBCKT OR4X8TS Y A B C D VSS VDD
X0 VDD nmin Y VDD LPPFET W=4.94U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=3.68U L=0.12U M=1 
X10 VDD D hnet14 VDD LPPFET W=1.18U L=0.12U M=1 
X11 hnet14 C hnet13 VDD LPPFET W=1.18U L=0.12U M=1 
X12 hnet13 B hnet15 VDD LPPFET W=1.18U L=0.12U M=1 
X13 hnet15 A nmin VDD LPPFET W=1.18U L=0.12U M=1 
X14 VDD D hnet24 VDD LPPFET W=1.18U L=0.12U M=1 
X15 hnet24 C hnet16 VDD LPPFET W=1.18U L=0.12U M=1 
X16 hnet16 B hnet19 VDD LPPFET W=1.18U L=0.12U M=1 
X17 hnet19 A nmin VDD LPPFET W=1.18U L=0.12U M=1 
X2 nmin D VSS VSS LPNFET W=1.24U L=0.12U M=1 
X3 nmin C VSS VSS LPNFET W=1.24U L=0.12U M=1 
X4 nmin B VSS VSS LPNFET W=1.24U L=0.12U M=1 
X5 nmin A VSS VSS LPNFET W=1.24U L=0.12U M=1 
X6 VDD D hnet26 VDD LPPFET W=1.18U L=0.12U M=1 
X7 hnet26 C hnet23 VDD LPPFET W=1.18U L=0.12U M=1 
X8 hnet23 B hnet18 VDD LPPFET W=1.18U L=0.12U M=1 
X9 hnet18 A nmin VDD LPPFET W=1.18U L=0.12U M=1 
.ENDS OR4X8TS 

**** 
*.SUBCKT OR4XLTS Y A B C D 
.SUBCKT OR4XLTS Y A B C D VSS VDD
X0 VDD nmin Y VDD LPPFET W=0.42U L=0.12U M=1 
X1 Y nmin VSS VSS LPNFET W=0.28U L=0.12U M=1 
X2 nmin D VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 nmin C VSS VSS LPNFET W=0.2U L=0.12U M=1 
X4 nmin B VSS VSS LPNFET W=0.2U L=0.12U M=1 
X5 nmin A VSS VSS LPNFET W=0.2U L=0.12U M=1 
X6 VDD D hnet15 VDD LPPFET W=0.42U L=0.12U M=1 
X7 hnet15 C hnet18 VDD LPPFET W=0.42U L=0.12U M=1 
X8 hnet18 B hnet14 VDD LPPFET W=0.42U L=0.12U M=1 
X9 hnet14 A nmin VDD LPPFET W=0.42U L=0.12U M=1 
.ENDS OR4XLTS 

**** 
*.SUBCKT RF1R1WX1TS RB RW RWN WB WW 
.SUBCKT RF1R1WX1TS RB RW RWN WB WW VSS VDD
X0 hnet12 WB VSS VSS LPNFET W=0.2U L=0.12U M=1 
X1 nmwrbl WW hnet12 VSS LPNFET W=0.2U L=0.12U M=1 
X10 hnet30 RWN RB VDD LPPFET W=0.64U L=0.12U M=1 
X11 VDD q hnet30 VDD LPPFET W=0.64U L=0.12U M=1 
X12 VDD WW nmwrwl VDD LPPFET W=0.36U L=0.12U M=1 
X13 nmwrwl WW VSS VSS LPNFET W=0.2U L=0.12U M=1 
X14 VDD nmwrbl q VDD LPPFET W=0.4U L=0.12U M=1 
X15 q nmwrbl VSS VSS LPNFET W=0.18U L=0.12U M=1 
X2 hnet14 nmwrwl nmwrbl VDD LPPFET W=0.38U L=0.12U M=1 
X3 VDD WB hnet14 VDD LPPFET W=0.38U L=0.12U M=1 
X4 hnet20 q VSS VSS LPNFET W=0.2U L=0.12U M=1 
X5 nmwrbl nmwrwl hnet20 VSS LPNFET W=0.2U L=0.12U M=1 
X6 hnet22 WW nmwrbl VDD LPPFET W=0.28U L=0.12U M=1 
X7 VDD q hnet22 VDD LPPFET W=0.28U L=0.12U M=1 
X8 hnet28 q VSS VSS LPNFET W=0.42U L=0.12U M=1 
X9 RB RW hnet28 VSS LPNFET W=0.42U L=0.12U M=1 
.ENDS RF1R1WX1TS 

**** 
*.SUBCKT RF2R1WX1TS R1B R2B R1W R2W WB WW 
.SUBCKT RF2R1WX1TS R1B R2B R1W R2W WB WW VSS VDD
X0 hnet15 q VSS VSS LPNFET W=0.88U L=0.12U M=1 
X1 R2B R2W hnet15 VSS LPNFET W=0.88U L=0.12U M=1 
X10 hnet33 WW nmwrbl VDD LPPFET W=0.28U L=0.12U M=1 
X11 VDD q hnet33 VDD LPPFET W=0.28U L=0.12U M=1 
X12 hnet39 q VSS VSS LPNFET W=0.88U L=0.12U M=1 
X13 R1B R1W hnet39 VSS LPNFET W=0.88U L=0.12U M=1 
X14 hnet41 nmrdwl1 R1B VDD LPPFET W=1.26U L=0.12U M=1 
X15 VDD q hnet41 VDD LPPFET W=1.26U L=0.12U M=1 
X16 VDD R2W nmrdwl2 VDD LPPFET W=0.3U L=0.12U M=1 
X17 nmrdwl2 R2W VSS VSS LPNFET W=0.22U L=0.12U M=1 
X18 VDD R1W nmrdwl1 VDD LPPFET W=0.3U L=0.12U M=1 
X19 nmrdwl1 R1W VSS VSS LPNFET W=0.22U L=0.12U M=1 
X2 hnet17 nmrdwl2 R2B VDD LPPFET W=1.28U L=0.12U M=1 
X20 VDD WW nmwrwl VDD LPPFET W=0.28U L=0.12U M=1 
X21 nmwrwl WW VSS VSS LPNFET W=0.2U L=0.12U M=1 
X22 VDD nmwrbl q VDD LPPFET W=1.12U L=0.12U M=1 
X23 q nmwrbl VSS VSS LPNFET W=0.78U L=0.12U M=1 
X3 VDD q hnet17 VDD LPPFET W=1.28U L=0.12U M=1 
X4 hnet23 WB VSS VSS LPNFET W=0.6U L=0.12U M=1 
X5 nmwrbl WW hnet23 VSS LPNFET W=0.6U L=0.12U M=1 
X6 hnet25 nmwrwl nmwrbl VDD LPPFET W=0.86U L=0.12U M=1 
X7 VDD WB hnet25 VDD LPPFET W=0.86U L=0.12U M=1 
X8 hnet31 q VSS VSS LPNFET W=0.2U L=0.12U M=1 
X9 nmwrbl nmwrwl hnet31 VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS RF2R1WX1TS 

**** 
*.SUBCKT RFRDX1TS BRB RB 
.SUBCKT RFRDX1TS BRB RB VSS VDD
X0 VDD BRB RB VDD LPPFET W=0.28U L=0.38U M=1 
X1 RB BRB VSS VSS LPNFET W=0.2U L=0.76U M=1 
X2 VDD RB BRB VDD LPPFET W=0.64U L=0.12U M=1 
X3 BRB RB VSS VSS LPNFET W=0.46U L=0.12U M=1 
.ENDS RFRDX1TS 

**** 
*.SUBCKT RFRDX2TS BRB RB 
.SUBCKT RFRDX2TS BRB RB VSS VDD
X0 VDD BRB RB VDD LPPFET W=0.28U L=0.38U M=1 
X1 RB BRB VSS VSS LPNFET W=0.2U L=0.76U M=1 
X2 VDD RB BRB VDD LPPFET W=1.28U L=0.12U M=1 
X3 BRB RB VSS VSS LPNFET W=0.92U L=0.12U M=1 
.ENDS RFRDX2TS 

**** 
*.SUBCKT RFRDX4TS BRB RB 
.SUBCKT RFRDX4TS BRB RB VSS VDD
X0 VDD BRB RB VDD LPPFET W=0.28U L=0.38U M=1 
X1 RB BRB VSS VSS LPNFET W=0.2U L=0.76U M=1 
X2 VDD RB BRB VDD LPPFET W=2.56U L=0.12U M=1 
X3 BRB RB VSS VSS LPNFET W=1.84U L=0.12U M=1 
.ENDS RFRDX4TS 

**** 
*.SUBCKT SDFFHQX1TS Q CK D SE SI 
.SUBCKT SDFFHQX1TS Q CK D SE SI VSS VDD
X0 VDD c hnet24 VDD LPPFET W=0.58U L=0.12U M=1 
X1 hnet24 nmsi pm VDD LPPFET W=0.58U L=0.12U M=1 
X10 net95 c m VSS LPNFET W=0.48U L=0.12U M=1 
X11 hnet30 SI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X12 nmsi SE hnet30 VSS LPNFET W=0.2U L=0.12U M=1 
X13 hnet32 nmse nmsi VDD LPPFET W=0.28U L=0.12U M=1 
X14 VDD SI hnet32 VDD LPPFET W=0.28U L=0.12U M=1 
X15 hnet36 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X16 pm c hnet36 VSS LPNFET W=0.2U L=0.12U M=1 
X17 hnet38 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X18 VDD m hnet38 VDD LPPFET W=0.28U L=0.12U M=1 
X19 hnet42 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 hnet28 cn VSS VSS LPNFET W=0.42U L=0.12U M=1 
X20 net95 cn hnet42 VSS LPNFET W=0.2U L=0.12U M=1 
X21 hnet44 c net95 VDD LPPFET W=0.28U L=0.12U M=1 
X22 VDD s hnet44 VDD LPPFET W=0.28U L=0.12U M=1 
X23 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X24 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X25 VDD D nmin VDD LPPFET W=0.38U L=0.12U M=1 
X26 nmin D VSS VSS LPNFET W=0.28U L=0.12U M=1 
X27 VDD pm m VDD LPPFET W=0.96U L=0.12U M=1 
X28 m pm VSS VSS LPNFET W=0.5U L=0.12U M=1 
X29 VDD net95 s VDD LPPFET W=0.28U L=0.12U M=1 
X3 pm nmsi hnet28 VSS LPNFET W=0.42U L=0.12U M=1 
X30 s net95 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X31 VDD net95 Q VDD LPPFET W=0.74U L=0.12U M=1 
X32 Q net95 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X33 VDD net110 c VDD LPPFET W=0.84U L=0.12U M=1 
X34 c net110 VSS VSS LPNFET W=0.3U L=0.12U M=1 
X35 VDD CK net110 VDD LPPFET W=0.28U L=0.12U M=1 
X36 net110 CK VSS VSS LPNFET W=0.28U L=0.12U M=1 
X4 net69 CK VDD VDD LPPFET W=0.7U L=0.12U M=1 
X5 cn c net69 VDD LPPFET W=0.52U L=0.12U M=1 
X6 nmsi SE nmin VDD LPPFET W=0.38U L=0.12U M=1 
X7 net95 cn m VDD LPPFET W=0.96U L=0.12U M=1 
X8 cn CK VSS VSS LPNFET W=0.2U L=0.12U M=1 
X9 nmsi nmse nmin VSS LPNFET W=0.28U L=0.12U M=1 
.ENDS SDFFHQX1TS 

**** 
*.SUBCKT SDFFHQX2TS Q CK D SE SI 
.SUBCKT SDFFHQX2TS Q CK D SE SI VSS VDD
X0 VDD c hnet24 VDD LPPFET W=1U L=0.12U M=1 
X1 hnet24 nmsi pm VDD LPPFET W=1U L=0.12U M=1 
X10 net95 c m VSS LPNFET W=0.82U L=0.12U M=1 
X11 hnet30 SI VSS VSS LPNFET W=0.24U L=0.12U M=1 
X12 nmsi SE hnet30 VSS LPNFET W=0.24U L=0.12U M=1 
X13 hnet32 nmse nmsi VDD LPPFET W=0.34U L=0.12U M=1 
X14 VDD SI hnet32 VDD LPPFET W=0.34U L=0.12U M=1 
X15 hnet36 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X16 pm c hnet36 VSS LPNFET W=0.2U L=0.12U M=1 
X17 hnet38 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X18 VDD m hnet38 VDD LPPFET W=0.28U L=0.12U M=1 
X19 hnet42 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 hnet28 cn VSS VSS LPNFET W=0.72U L=0.12U M=1 
X20 net95 cn hnet42 VSS LPNFET W=0.2U L=0.12U M=1 
X21 hnet44 c net95 VDD LPPFET W=0.28U L=0.12U M=1 
X22 VDD s hnet44 VDD LPPFET W=0.28U L=0.12U M=1 
X23 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X24 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X25 VDD D nmin VDD LPPFET W=0.68U L=0.12U M=1 
X26 nmin D VSS VSS LPNFET W=0.5U L=0.12U M=1 
X27 VDD pm m VDD LPPFET W=1.64U L=0.12U M=1 
X28 m pm VSS VSS LPNFET W=0.86U L=0.12U M=1 
X29 VDD net95 s VDD LPPFET W=0.28U L=0.12U M=1 
X3 pm nmsi hnet28 VSS LPNFET W=0.72U L=0.12U M=1 
X30 s net95 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X31 VDD net95 Q VDD LPPFET W=1.3U L=0.12U M=1 
X32 Q net95 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X33 VDD net110 c VDD LPPFET W=1.18U L=0.12U M=1 
X34 c net110 VSS VSS LPNFET W=0.42U L=0.12U M=1 
X35 VDD CK net110 VDD LPPFET W=0.32U L=0.12U M=1 
X36 net110 CK VSS VSS LPNFET W=0.32U L=0.12U M=1 
X4 net67 CK VDD VDD LPPFET W=0.9U L=0.12U M=1 
X5 cn c net67 VDD LPPFET W=0.68U L=0.12U M=1 
X6 nmsi SE nmin VDD LPPFET W=0.68U L=0.12U M=1 
X7 net95 cn m VDD LPPFET W=1.64U L=0.12U M=1 
X8 cn CK VSS VSS LPNFET W=0.26U L=0.12U M=1 
X9 nmsi nmse nmin VSS LPNFET W=0.5U L=0.12U M=1 
.ENDS SDFFHQX2TS 

**** 
*.SUBCKT SDFFHQX4TS Q CK D SE SI 
.SUBCKT SDFFHQX4TS Q CK D SE SI VSS VDD
X0 hnet26 cn VSS VSS LPNFET W=0.6U L=0.12U M=1 
X1 pm nmsi hnet26 VSS LPNFET W=0.6U L=0.12U M=1 
X10 net75 CK VDD VDD LPPFET W=0.84U L=0.12U M=1 
X11 cn c net75 VDD LPPFET W=0.64U L=0.12U M=1 
X12 nmsi SE nmin VDD LPPFET W=1.22U L=0.12U M=1 
X13 net101 cn m VDD LPPFET W=3U L=0.12U M=1 
X14 cn CK VSS VSS LPNFET W=0.48U L=0.12U M=1 
X15 nmsi nmse nmin VSS LPNFET W=0.88U L=0.12U M=1 
X16 net101 c m VSS LPNFET W=1.5U L=0.12U M=1 
X17 hnet33 SI VSS VSS LPNFET W=0.44U L=0.12U M=1 
X18 nmsi SE hnet33 VSS LPNFET W=0.44U L=0.12U M=1 
X19 hnet35 nmse nmsi VDD LPPFET W=0.62U L=0.12U M=1 
X2 hnet22 cn VSS VSS LPNFET W=0.6U L=0.12U M=1 
X20 VDD SI hnet35 VDD LPPFET W=0.62U L=0.12U M=1 
X21 hnet39 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X22 pm c hnet39 VSS LPNFET W=0.2U L=0.12U M=1 
X23 hnet41 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X24 VDD m hnet41 VDD LPPFET W=0.28U L=0.12U M=1 
X25 hnet45 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X26 net101 cn hnet45 VSS LPNFET W=0.2U L=0.12U M=1 
X27 hnet47 c net101 VDD LPPFET W=0.28U L=0.12U M=1 
X28 VDD s hnet47 VDD LPPFET W=0.28U L=0.12U M=1 
X29 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X3 pm nmsi hnet22 VSS LPNFET W=0.6U L=0.12U M=1 
X30 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X31 VDD D nmin VDD LPPFET W=1.22U L=0.12U M=1 
X32 nmin D VSS VSS LPNFET W=0.88U L=0.12U M=1 
X33 VDD pm m VDD LPPFET W=2.6U L=0.12U M=1 
X34 m pm VSS VSS LPNFET W=1.56U L=0.12U M=1 
X35 VDD net101 s VDD LPPFET W=0.28U L=0.12U M=1 
X36 s net101 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X37 VDD net101 Q VDD LPPFET W=2.62U L=0.12U M=1 
X38 Q net101 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X39 VDD net116 c VDD LPPFET W=2U L=0.12U M=1 
X4 VDD c hnet31 VDD LPPFET W=0.9U L=0.12U M=1 
X40 c net116 VSS VSS LPNFET W=0.72U L=0.12U M=1 
X41 VDD CK net116 VDD LPPFET W=0.54U L=0.12U M=1 
X42 net116 CK VSS VSS LPNFET W=0.54U L=0.12U M=1 
X5 hnet31 nmsi pm VDD LPPFET W=0.9U L=0.12U M=1 
X6 VDD c hnet28 VDD LPPFET W=0.9U L=0.12U M=1 
X7 hnet28 nmsi pm VDD LPPFET W=0.9U L=0.12U M=1 
X8 cn c net70 VDD LPPFET W=0.64U L=0.12U M=1 
X9 net70 CK VDD VDD LPPFET W=0.84U L=0.12U M=1 
.ENDS SDFFHQX4TS 

**** 
*.SUBCKT SDFFHQX8TS Q CK D SE SI 
.SUBCKT SDFFHQX8TS Q CK D SE SI VSS VDD
X0 hnet26 cn VSS VSS LPNFET W=0.6U L=0.12U M=1 
X1 pm nmsi hnet26 VSS LPNFET W=0.6U L=0.12U M=1 
X10 net75 CK VDD VDD LPPFET W=0.84U L=0.12U M=1 
X11 cn c net75 VDD LPPFET W=0.64U L=0.12U M=1 
X12 nmsi SE nmin VDD LPPFET W=1.22U L=0.12U M=1 
X13 net101 cn m VDD LPPFET W=3U L=0.12U M=1 
X14 cn CK VSS VSS LPNFET W=0.48U L=0.12U M=1 
X15 nmsi nmse nmin VSS LPNFET W=0.88U L=0.12U M=1 
X16 net101 c m VSS LPNFET W=1.5U L=0.12U M=1 
X17 hnet33 SI VSS VSS LPNFET W=0.44U L=0.12U M=1 
X18 nmsi SE hnet33 VSS LPNFET W=0.44U L=0.12U M=1 
X19 hnet35 nmse nmsi VDD LPPFET W=0.62U L=0.12U M=1 
X2 hnet22 cn VSS VSS LPNFET W=0.6U L=0.12U M=1 
X20 VDD SI hnet35 VDD LPPFET W=0.62U L=0.12U M=1 
X21 hnet39 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X22 pm c hnet39 VSS LPNFET W=0.2U L=0.12U M=1 
X23 hnet41 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X24 VDD m hnet41 VDD LPPFET W=0.28U L=0.12U M=1 
X25 hnet45 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X26 net101 cn hnet45 VSS LPNFET W=0.2U L=0.12U M=1 
X27 hnet47 c net101 VDD LPPFET W=0.28U L=0.12U M=1 
X28 VDD s hnet47 VDD LPPFET W=0.28U L=0.12U M=1 
X29 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X3 pm nmsi hnet22 VSS LPNFET W=0.6U L=0.12U M=1 
X30 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X31 VDD D nmin VDD LPPFET W=1.22U L=0.12U M=1 
X32 nmin D VSS VSS LPNFET W=0.88U L=0.12U M=1 
X33 VDD pm m VDD LPPFET W=2.6U L=0.12U M=1 
X34 m pm VSS VSS LPNFET W=1.56U L=0.12U M=1 
X35 VDD net101 s VDD LPPFET W=0.28U L=0.12U M=1 
X36 s net101 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X37 VDD net101 Q VDD LPPFET W=5.2U L=0.12U M=1 
X38 Q net101 VSS VSS LPNFET W=3.68U L=0.12U M=1 
X39 VDD net116 c VDD LPPFET W=2U L=0.12U M=1 
X4 VDD c hnet31 VDD LPPFET W=0.9U L=0.12U M=1 
X40 c net116 VSS VSS LPNFET W=0.72U L=0.12U M=1 
X41 VDD CK net116 VDD LPPFET W=0.54U L=0.12U M=1 
X42 net116 CK VSS VSS LPNFET W=0.54U L=0.12U M=1 
X5 hnet31 nmsi pm VDD LPPFET W=0.9U L=0.12U M=1 
X6 VDD c hnet28 VDD LPPFET W=0.9U L=0.12U M=1 
X7 hnet28 nmsi pm VDD LPPFET W=0.9U L=0.12U M=1 
X8 cn c net70 VDD LPPFET W=0.64U L=0.12U M=1 
X9 net70 CK VDD VDD LPPFET W=0.84U L=0.12U M=1 
.ENDS SDFFHQX8TS 

**** 
*.SUBCKT SDFFNSRX1TS Q QN CKN D RN SE SI SN 
.SUBCKT SDFFNSRX1TS Q QN CKN D RN SE SI SN VSS VDD
X0 VDD D hnet32 VDD LPPFET W=0.28U L=0.12U M=1 
X1 hnet32 SE nminsi VDD LPPFET W=0.28U L=0.12U M=1 
X10 net148 c net106 VDD LPPFET W=0.28U L=0.12U M=1 
X11 net148 cn m VDD LPPFET W=0.28U L=0.12U M=1 
X12 net117 D VSS VSS LPNFET W=0.2U L=0.12U M=1 
X13 nminsi nmse net117 VSS LPNFET W=0.2U L=0.12U M=1 
X14 net121 SI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X15 nminsi SE net121 VSS LPNFET W=0.2U L=0.12U M=1 
X16 pm cn nminsi VSS LPNFET W=0.2U L=0.12U M=1 
X17 m net159 net142 VSS LPNFET W=0.2U L=0.12U M=1 
X18 m pm net142 VSS LPNFET W=0.3U L=0.12U M=1 
X19 net148 net159 net142 VSS LPNFET W=0.2U L=0.12U M=1 
X2 VDD SI hnet36 VDD LPPFET W=0.28U L=0.12U M=1 
X20 net139 s net142 VSS LPNFET W=0.2U L=0.12U M=1 
X21 net142 SN VSS VSS LPNFET W=0.4U L=0.12U M=1 
X22 net148 cn net139 VSS LPNFET W=0.2U L=0.12U M=1 
X23 net148 c m VSS LPNFET W=0.2U L=0.12U M=1 
X24 hnet38 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X25 pm c hnet38 VSS LPNFET W=0.2U L=0.12U M=1 
X26 hnet40 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X27 VDD m hnet40 VDD LPPFET W=0.28U L=0.12U M=1 
X28 VDD s net153 VDD LPPFET W=0.28U L=0.12U M=1 
X29 net153 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 hnet36 nmse nminsi VDD LPPFET W=0.28U L=0.12U M=1 
X30 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X31 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X32 VDD s Q VDD LPPFET W=0.64U L=0.12U M=1 
X33 Q s VSS VSS LPNFET W=0.46U L=0.12U M=1 
X34 VDD RN net159 VDD LPPFET W=0.28U L=0.12U M=1 
X35 net159 RN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X36 VDD net148 s VDD LPPFET W=0.28U L=0.12U M=1 
X37 s net148 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X38 VDD net153 QN VDD LPPFET W=0.64U L=0.12U M=1 
X39 QN net153 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X4 pm c nminsi VDD LPPFET W=0.28U L=0.12U M=1 
X40 VDD CKN c VDD LPPFET W=0.42U L=0.12U M=1 
X41 c CKN VSS VSS LPNFET W=0.3U L=0.12U M=1 
X42 VDD c cn VDD LPPFET W=0.28U L=0.12U M=1 
X43 cn c VSS VSS LPNFET W=0.2U L=0.12U M=1 
X5 m SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X6 m pm net96 VDD LPPFET W=0.42U L=0.12U M=1 
X7 net96 net159 VDD VDD LPPFET W=0.56U L=0.12U M=1 
X8 net148 SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X9 net106 s net96 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS SDFFNSRX1TS 

**** 
*.SUBCKT SDFFNSRX2TS Q QN CKN D RN SE SI SN 
.SUBCKT SDFFNSRX2TS Q QN CKN D RN SE SI SN VSS VDD
X0 VDD D hnet32 VDD LPPFET W=0.28U L=0.12U M=1 
X1 hnet32 SE nminsi VDD LPPFET W=0.28U L=0.12U M=1 
X10 net148 c net106 VDD LPPFET W=0.28U L=0.12U M=1 
X11 net148 cn m VDD LPPFET W=0.28U L=0.12U M=1 
X12 net117 D VSS VSS LPNFET W=0.2U L=0.12U M=1 
X13 nminsi nmse net117 VSS LPNFET W=0.2U L=0.12U M=1 
X14 net123 SI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X15 nminsi SE net123 VSS LPNFET W=0.2U L=0.12U M=1 
X16 pm cn nminsi VSS LPNFET W=0.2U L=0.12U M=1 
X17 m net159 net142 VSS LPNFET W=0.2U L=0.12U M=1 
X18 m pm net142 VSS LPNFET W=0.3U L=0.12U M=1 
X19 net148 net159 net142 VSS LPNFET W=0.2U L=0.12U M=1 
X2 VDD SI hnet36 VDD LPPFET W=0.28U L=0.12U M=1 
X20 net144 s net142 VSS LPNFET W=0.2U L=0.12U M=1 
X21 net142 SN VSS VSS LPNFET W=0.4U L=0.12U M=1 
X22 net148 cn net144 VSS LPNFET W=0.2U L=0.12U M=1 
X23 net148 c m VSS LPNFET W=0.2U L=0.12U M=1 
X24 hnet38 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X25 pm c hnet38 VSS LPNFET W=0.2U L=0.12U M=1 
X26 hnet40 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X27 VDD m hnet40 VDD LPPFET W=0.28U L=0.12U M=1 
X28 VDD s net153 VDD LPPFET W=0.3U L=0.12U M=1 
X29 net153 s VSS VSS LPNFET W=0.22U L=0.12U M=1 
X3 hnet36 nmse nminsi VDD LPPFET W=0.28U L=0.12U M=1 
X30 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X31 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X32 VDD s Q VDD LPPFET W=1.28U L=0.12U M=1 
X33 Q s VSS VSS LPNFET W=0.92U L=0.12U M=1 
X34 VDD RN net159 VDD LPPFET W=0.28U L=0.12U M=1 
X35 net159 RN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X36 VDD net148 s VDD LPPFET W=0.34U L=0.12U M=1 
X37 s net148 VSS VSS LPNFET W=0.26U L=0.12U M=1 
X38 VDD net153 QN VDD LPPFET W=1.28U L=0.12U M=1 
X39 QN net153 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X4 pm c nminsi VDD LPPFET W=0.28U L=0.12U M=1 
X40 VDD CKN c VDD LPPFET W=0.42U L=0.12U M=1 
X41 c CKN VSS VSS LPNFET W=0.3U L=0.12U M=1 
X42 VDD c cn VDD LPPFET W=0.28U L=0.12U M=1 
X43 cn c VSS VSS LPNFET W=0.2U L=0.12U M=1 
X5 m SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X6 m pm net96 VDD LPPFET W=0.42U L=0.12U M=1 
X7 net96 net159 VDD VDD LPPFET W=0.56U L=0.12U M=1 
X8 net148 SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X9 net106 s net96 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS SDFFNSRX2TS 

**** 
*.SUBCKT SDFFNSRX4TS Q QN CKN D RN SE SI SN 
.SUBCKT SDFFNSRX4TS Q QN CKN D RN SE SI SN VSS VDD
X0 VDD D hnet32 VDD LPPFET W=0.28U L=0.12U M=1 
X1 hnet32 SE nminsi VDD LPPFET W=0.28U L=0.12U M=1 
X10 net148 c net106 VDD LPPFET W=0.28U L=0.12U M=1 
X11 net148 cn m VDD LPPFET W=0.3U L=0.12U M=1 
X12 net117 D VSS VSS LPNFET W=0.2U L=0.12U M=1 
X13 nminsi nmse net117 VSS LPNFET W=0.2U L=0.12U M=1 
X14 net123 SI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X15 nminsi SE net123 VSS LPNFET W=0.2U L=0.12U M=1 
X16 pm cn nminsi VSS LPNFET W=0.2U L=0.12U M=1 
X17 m net159 net142 VSS LPNFET W=0.2U L=0.12U M=1 
X18 m pm net142 VSS LPNFET W=0.34U L=0.12U M=1 
X19 net148 net159 net142 VSS LPNFET W=0.2U L=0.12U M=1 
X2 VDD SI hnet36 VDD LPPFET W=0.28U L=0.12U M=1 
X20 net144 s net142 VSS LPNFET W=0.2U L=0.12U M=1 
X21 net142 SN VSS VSS LPNFET W=0.46U L=0.12U M=1 
X22 net148 cn net144 VSS LPNFET W=0.2U L=0.12U M=1 
X23 net148 c m VSS LPNFET W=0.22U L=0.12U M=1 
X24 hnet38 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X25 pm c hnet38 VSS LPNFET W=0.2U L=0.12U M=1 
X26 hnet40 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X27 VDD m hnet40 VDD LPPFET W=0.28U L=0.12U M=1 
X28 VDD s net153 VDD LPPFET W=0.62U L=0.12U M=1 
X29 net153 s VSS VSS LPNFET W=0.4U L=0.12U M=1 
X3 hnet36 nmse nminsi VDD LPPFET W=0.28U L=0.12U M=1 
X30 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X31 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X32 VDD s Q VDD LPPFET W=2.4U L=0.12U M=1 
X33 Q s VSS VSS LPNFET W=1.84U L=0.12U M=1 
X34 VDD RN net159 VDD LPPFET W=0.28U L=0.12U M=1 
X35 net159 RN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X36 VDD net148 s VDD LPPFET W=0.66U L=0.12U M=1 
X37 s net148 VSS VSS LPNFET W=0.44U L=0.12U M=1 
X38 VDD net153 QN VDD LPPFET W=2.4U L=0.12U M=1 
X39 QN net153 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X4 pm c nminsi VDD LPPFET W=0.28U L=0.12U M=1 
X40 VDD CKN c VDD LPPFET W=0.44U L=0.12U M=1 
X41 c CKN VSS VSS LPNFET W=0.32U L=0.12U M=1 
X42 VDD c cn VDD LPPFET W=0.28U L=0.12U M=1 
X43 cn c VSS VSS LPNFET W=0.2U L=0.12U M=1 
X5 m SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X6 m pm net96 VDD LPPFET W=0.46U L=0.12U M=1 
X7 net96 net159 VDD VDD LPPFET W=0.62U L=0.12U M=1 
X8 net148 SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X9 net106 s net96 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS SDFFNSRX4TS 

**** 
*.SUBCKT SDFFNSRXLTS Q QN CKN D RN SE SI SN 
.SUBCKT SDFFNSRXLTS Q QN CKN D RN SE SI SN VSS VDD
X0 VDD D hnet32 VDD LPPFET W=0.28U L=0.12U M=1 
X1 hnet32 SE nminsi VDD LPPFET W=0.28U L=0.12U M=1 
X10 net148 c net106 VDD LPPFET W=0.28U L=0.12U M=1 
X11 net148 cn m VDD LPPFET W=0.28U L=0.12U M=1 
X12 net117 D VSS VSS LPNFET W=0.2U L=0.12U M=1 
X13 nminsi nmse net117 VSS LPNFET W=0.2U L=0.12U M=1 
X14 net123 SI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X15 nminsi SE net123 VSS LPNFET W=0.2U L=0.12U M=1 
X16 pm cn nminsi VSS LPNFET W=0.2U L=0.12U M=1 
X17 m net159 net142 VSS LPNFET W=0.2U L=0.12U M=1 
X18 m pm net142 VSS LPNFET W=0.3U L=0.12U M=1 
X19 net148 net159 net142 VSS LPNFET W=0.2U L=0.12U M=1 
X2 VDD SI hnet36 VDD LPPFET W=0.28U L=0.12U M=1 
X20 net144 s net142 VSS LPNFET W=0.2U L=0.12U M=1 
X21 net142 SN VSS VSS LPNFET W=0.4U L=0.12U M=1 
X22 net148 cn net144 VSS LPNFET W=0.2U L=0.12U M=1 
X23 net148 c m VSS LPNFET W=0.2U L=0.12U M=1 
X24 hnet38 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X25 pm c hnet38 VSS LPNFET W=0.2U L=0.12U M=1 
X26 hnet40 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X27 VDD m hnet40 VDD LPPFET W=0.28U L=0.12U M=1 
X28 VDD s net153 VDD LPPFET W=0.28U L=0.12U M=1 
X29 net153 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 hnet36 nmse nminsi VDD LPPFET W=0.28U L=0.12U M=1 
X30 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X31 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X32 VDD s Q VDD LPPFET W=0.34U L=0.12U M=1 
X33 Q s VSS VSS LPNFET W=0.24U L=0.12U M=1 
X34 VDD RN net159 VDD LPPFET W=0.28U L=0.12U M=1 
X35 net159 RN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X36 VDD net148 s VDD LPPFET W=0.28U L=0.12U M=1 
X37 s net148 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X38 VDD net153 QN VDD LPPFET W=0.34U L=0.12U M=1 
X39 QN net153 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X4 pm c nminsi VDD LPPFET W=0.28U L=0.12U M=1 
X40 VDD CKN c VDD LPPFET W=0.42U L=0.12U M=1 
X41 c CKN VSS VSS LPNFET W=0.3U L=0.12U M=1 
X42 VDD c cn VDD LPPFET W=0.28U L=0.12U M=1 
X43 cn c VSS VSS LPNFET W=0.2U L=0.12U M=1 
X5 m SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X6 m pm net96 VDD LPPFET W=0.42U L=0.12U M=1 
X7 net96 net159 VDD VDD LPPFET W=0.56U L=0.12U M=1 
X8 net148 SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X9 net106 s net96 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS SDFFNSRXLTS 

**** 
*.SUBCKT SDFFQX1TS Q CK D SE SI 
.SUBCKT SDFFQX1TS Q CK D SE SI VSS VDD
X0 net56 SE net65 VSS LPNFET W=0.2U L=0.12U M=1 
X1 net56 D net59 VSS LPNFET W=0.2U L=0.12U M=1 
X10 net83 SI VDD VDD LPPFET W=0.28U L=0.12U M=1 
X11 net68 cn m VDD LPPFET W=0.28U L=0.12U M=1 
X12 hnet24 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X13 net68 cn hnet24 VSS LPNFET W=0.2U L=0.12U M=1 
X14 hnet26 c net68 VDD LPPFET W=0.28U L=0.12U M=1 
X15 VDD s hnet26 VDD LPPFET W=0.28U L=0.12U M=1 
X16 hnet30 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X17 pm c hnet30 VSS LPNFET W=0.2U L=0.12U M=1 
X18 hnet32 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X19 VDD m hnet32 VDD LPPFET W=0.28U L=0.12U M=1 
X2 net59 nmse VSS VSS LPNFET W=0.2U L=0.12U M=1 
X20 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X21 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X22 VDD net68 s VDD LPPFET W=0.28U L=0.12U M=1 
X23 s net68 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X24 VDD pm m VDD LPPFET W=0.28U L=0.12U M=1 
X25 m pm VSS VSS LPNFET W=0.2U L=0.12U M=1 
X26 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X27 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X28 VDD CK cn VDD LPPFET W=0.38U L=0.12U M=1 
X29 cn CK VSS VSS LPNFET W=0.28U L=0.12U M=1 
X3 pm cn net56 VSS LPNFET W=0.2U L=0.12U M=1 
X30 VDD s Q VDD LPPFET W=0.64U L=0.12U M=1 
X31 Q s VSS VSS LPNFET W=0.48U L=0.12U M=1 
X4 net65 SI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X5 net68 c m VSS LPNFET W=0.2U L=0.12U M=1 
X6 net71 D net74 VDD LPPFET W=0.28U L=0.12U M=1 
X7 net74 SE VDD VDD LPPFET W=0.28U L=0.12U M=1 
X8 net71 nmse net83 VDD LPPFET W=0.28U L=0.12U M=1 
X9 pm c net71 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS SDFFQX1TS 

**** 
*.SUBCKT SDFFQX2TS Q CK D SE SI 
.SUBCKT SDFFQX2TS Q CK D SE SI VSS VDD
X0 net56 SE net65 VSS LPNFET W=0.2U L=0.12U M=1 
X1 net56 D net59 VSS LPNFET W=0.2U L=0.12U M=1 
X10 net83 SI VDD VDD LPPFET W=0.28U L=0.12U M=1 
X11 net68 cn m VDD LPPFET W=0.28U L=0.12U M=1 
X12 hnet24 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X13 net68 cn hnet24 VSS LPNFET W=0.2U L=0.12U M=1 
X14 hnet26 c net68 VDD LPPFET W=0.28U L=0.12U M=1 
X15 VDD s hnet26 VDD LPPFET W=0.28U L=0.12U M=1 
X16 hnet30 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X17 pm c hnet30 VSS LPNFET W=0.2U L=0.12U M=1 
X18 hnet32 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X19 VDD m hnet32 VDD LPPFET W=0.28U L=0.12U M=1 
X2 net59 nmse VSS VSS LPNFET W=0.2U L=0.12U M=1 
X20 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X21 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X22 VDD net68 s VDD LPPFET W=0.28U L=0.12U M=1 
X23 s net68 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X24 VDD pm m VDD LPPFET W=0.28U L=0.12U M=1 
X25 m pm VSS VSS LPNFET W=0.2U L=0.12U M=1 
X26 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X27 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X28 VDD CK cn VDD LPPFET W=0.38U L=0.12U M=1 
X29 cn CK VSS VSS LPNFET W=0.28U L=0.12U M=1 
X3 pm cn net56 VSS LPNFET W=0.2U L=0.12U M=1 
X30 VDD s Q VDD LPPFET W=1.28U L=0.12U M=1 
X31 Q s VSS VSS LPNFET W=0.92U L=0.12U M=1 
X4 net65 SI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X5 net68 c m VSS LPNFET W=0.2U L=0.12U M=1 
X6 net71 D net74 VDD LPPFET W=0.28U L=0.12U M=1 
X7 net74 SE VDD VDD LPPFET W=0.28U L=0.12U M=1 
X8 net71 nmse net83 VDD LPPFET W=0.28U L=0.12U M=1 
X9 pm c net71 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS SDFFQX2TS 

**** 
*.SUBCKT SDFFQX4TS Q CK D SE SI 
.SUBCKT SDFFQX4TS Q CK D SE SI VSS VDD
X0 net56 SE net65 VSS LPNFET W=0.2U L=0.12U M=1 
X1 net56 D net59 VSS LPNFET W=0.2U L=0.12U M=1 
X10 net83 SI VDD VDD LPPFET W=0.28U L=0.12U M=1 
X11 net68 cn m VDD LPPFET W=0.28U L=0.12U M=1 
X12 hnet24 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X13 net68 cn hnet24 VSS LPNFET W=0.2U L=0.12U M=1 
X14 hnet26 c net68 VDD LPPFET W=0.28U L=0.12U M=1 
X15 VDD s hnet26 VDD LPPFET W=0.28U L=0.12U M=1 
X16 hnet30 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X17 pm c hnet30 VSS LPNFET W=0.2U L=0.12U M=1 
X18 hnet32 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X19 VDD m hnet32 VDD LPPFET W=0.28U L=0.12U M=1 
X2 net59 nmse VSS VSS LPNFET W=0.2U L=0.12U M=1 
X20 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X21 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X22 VDD net68 s VDD LPPFET W=0.5U L=0.12U M=1 
X23 s net68 VSS VSS LPNFET W=0.36U L=0.12U M=1 
X24 VDD pm m VDD LPPFET W=0.28U L=0.12U M=1 
X25 m pm VSS VSS LPNFET W=0.2U L=0.12U M=1 
X26 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X27 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X28 VDD CK cn VDD LPPFET W=0.38U L=0.12U M=1 
X29 cn CK VSS VSS LPNFET W=0.28U L=0.12U M=1 
X3 pm cn net56 VSS LPNFET W=0.2U L=0.12U M=1 
X30 VDD s Q VDD LPPFET W=2.56U L=0.12U M=1 
X31 Q s VSS VSS LPNFET W=1.84U L=0.12U M=1 
X4 net65 SI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X5 net68 c m VSS LPNFET W=0.2U L=0.12U M=1 
X6 net71 D net74 VDD LPPFET W=0.28U L=0.12U M=1 
X7 net74 SE VDD VDD LPPFET W=0.28U L=0.12U M=1 
X8 net71 nmse net83 VDD LPPFET W=0.28U L=0.12U M=1 
X9 pm c net71 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS SDFFQX4TS 

**** 
*.SUBCKT SDFFQXLTS Q CK D SE SI 
.SUBCKT SDFFQXLTS Q CK D SE SI VSS VDD
X0 net56 SE net65 VSS LPNFET W=0.2U L=0.12U M=1 
X1 net56 D net59 VSS LPNFET W=0.2U L=0.12U M=1 
X10 net83 SI VDD VDD LPPFET W=0.28U L=0.12U M=1 
X11 net68 cn m VDD LPPFET W=0.28U L=0.12U M=1 
X12 hnet24 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X13 net68 cn hnet24 VSS LPNFET W=0.2U L=0.12U M=1 
X14 hnet26 c net68 VDD LPPFET W=0.28U L=0.12U M=1 
X15 VDD s hnet26 VDD LPPFET W=0.28U L=0.12U M=1 
X16 hnet30 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X17 pm c hnet30 VSS LPNFET W=0.2U L=0.12U M=1 
X18 hnet32 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X19 VDD m hnet32 VDD LPPFET W=0.28U L=0.12U M=1 
X2 net59 nmse VSS VSS LPNFET W=0.2U L=0.12U M=1 
X20 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X21 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X22 VDD net68 s VDD LPPFET W=0.28U L=0.12U M=1 
X23 s net68 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X24 VDD pm m VDD LPPFET W=0.28U L=0.12U M=1 
X25 m pm VSS VSS LPNFET W=0.2U L=0.12U M=1 
X26 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X27 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X28 VDD CK cn VDD LPPFET W=0.38U L=0.12U M=1 
X29 cn CK VSS VSS LPNFET W=0.28U L=0.12U M=1 
X3 pm cn net56 VSS LPNFET W=0.2U L=0.12U M=1 
X30 VDD s Q VDD LPPFET W=0.34U L=0.12U M=1 
X31 Q s VSS VSS LPNFET W=0.24U L=0.12U M=1 
X4 net65 SI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X5 net68 c m VSS LPNFET W=0.2U L=0.12U M=1 
X6 net71 D net74 VDD LPPFET W=0.28U L=0.12U M=1 
X7 net74 SE VDD VDD LPPFET W=0.28U L=0.12U M=1 
X8 net71 nmse net83 VDD LPPFET W=0.28U L=0.12U M=1 
X9 pm c net71 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS SDFFQXLTS 

**** 
*.SUBCKT SDFFRHQX1TS Q CK D RN SE SI 
.SUBCKT SDFFRHQX1TS Q CK D RN SE SI VSS VDD
X0 VDD c hnet28 VDD LPPFET W=0.62U L=0.12U M=1 
X1 hnet28 nmsi pm VDD LPPFET W=0.62U L=0.12U M=1 
X10 net122 c net91 VDD LPPFET W=0.28U L=0.12U M=1 
X11 net91 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X12 m RN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X13 m pm VDD VDD LPPFET W=0.96U L=0.12U M=1 
X14 net122 cn m VDD LPPFET W=0.92U L=0.12U M=1 
X15 cn CK VSS VSS LPNFET W=0.2U L=0.12U M=1 
X16 nmsi nmse nmin VSS LPNFET W=0.3U L=0.12U M=1 
X17 net115 RN net112 VSS LPNFET W=0.2U L=0.12U M=1 
X18 net122 cn net115 VSS LPNFET W=0.2U L=0.12U M=1 
X19 net112 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 hnet32 cn VSS VSS LPNFET W=0.44U L=0.12U M=1 
X20 net122 c m VSS LPNFET W=0.48U L=0.12U M=1 
X21 hnet38 SI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X22 nmsi SE hnet38 VSS LPNFET W=0.2U L=0.12U M=1 
X23 hnet40 nmse nmsi VDD LPPFET W=0.28U L=0.12U M=1 
X24 VDD SI hnet40 VDD LPPFET W=0.28U L=0.12U M=1 
X25 hnet44 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X26 pm c hnet44 VSS LPNFET W=0.2U L=0.12U M=1 
X27 hnet46 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X28 VDD m hnet46 VDD LPPFET W=0.28U L=0.12U M=1 
X29 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X3 pm nmsi hnet32 VSS LPNFET W=0.44U L=0.12U M=1 
X30 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X31 VDD D nmin VDD LPPFET W=0.42U L=0.12U M=1 
X32 nmin D VSS VSS LPNFET W=0.3U L=0.12U M=1 
X33 VDD net122 s VDD LPPFET W=0.28U L=0.12U M=1 
X34 s net122 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X35 VDD net122 Q VDD LPPFET W=0.74U L=0.12U M=1 
X36 Q net122 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X37 VDD net141 c VDD LPPFET W=0.84U L=0.12U M=1 
X38 c net141 VSS VSS LPNFET W=0.3U L=0.12U M=1 
X39 VDD CK net141 VDD LPPFET W=0.28U L=0.12U M=1 
X4 hnet36 RN VSS VSS LPNFET W=0.58U L=0.12U M=1 
X40 net141 CK VSS VSS LPNFET W=0.28U L=0.12U M=1 
X5 m pm hnet36 VSS LPNFET W=0.58U L=0.12U M=1 
X6 net80 CK VDD VDD LPPFET W=0.7U L=0.12U M=1 
X7 cn c net80 VDD LPPFET W=0.52U L=0.12U M=1 
X8 nmsi SE nmin VDD LPPFET W=0.42U L=0.12U M=1 
X9 net122 RN VDD VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS SDFFRHQX1TS 

**** 
*.SUBCKT SDFFRHQX2TS Q CK D RN SE SI 
.SUBCKT SDFFRHQX2TS Q CK D RN SE SI VSS VDD
X0 VDD c hnet28 VDD LPPFET W=1.02U L=0.12U M=1 
X1 hnet28 nmsi pm VDD LPPFET W=1.02U L=0.12U M=1 
X10 net122 c net91 VDD LPPFET W=0.28U L=0.12U M=1 
X11 net91 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X12 m RN VDD VDD LPPFET W=0.4U L=0.12U M=1 
X13 m pm VDD VDD LPPFET W=1.64U L=0.12U M=1 
X14 net122 cn m VDD LPPFET W=1.64U L=0.12U M=1 
X15 cn CK VSS VSS LPNFET W=0.28U L=0.12U M=1 
X16 nmsi nmse nmin VSS LPNFET W=0.5U L=0.12U M=1 
X17 net115 RN net112 VSS LPNFET W=0.2U L=0.12U M=1 
X18 net122 cn net115 VSS LPNFET W=0.2U L=0.12U M=1 
X19 net112 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 hnet32 cn VSS VSS LPNFET W=0.74U L=0.12U M=1 
X20 net122 c m VSS LPNFET W=0.74U L=0.12U M=1 
X21 hnet38 SI VSS VSS LPNFET W=0.28U L=0.12U M=1 
X22 nmsi SE hnet38 VSS LPNFET W=0.28U L=0.12U M=1 
X23 hnet40 nmse nmsi VDD LPPFET W=0.36U L=0.12U M=1 
X24 VDD SI hnet40 VDD LPPFET W=0.36U L=0.12U M=1 
X25 hnet44 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X26 pm c hnet44 VSS LPNFET W=0.2U L=0.12U M=1 
X27 hnet46 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X28 VDD m hnet46 VDD LPPFET W=0.28U L=0.12U M=1 
X29 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X3 pm nmsi hnet32 VSS LPNFET W=0.74U L=0.12U M=1 
X30 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X31 VDD D nmin VDD LPPFET W=0.7U L=0.12U M=1 
X32 nmin D VSS VSS LPNFET W=0.5U L=0.12U M=1 
X33 VDD net122 s VDD LPPFET W=0.28U L=0.12U M=1 
X34 s net122 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X35 VDD net122 Q VDD LPPFET W=1.3U L=0.12U M=1 
X36 Q net122 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X37 VDD net141 c VDD LPPFET W=1.16U L=0.12U M=1 
X38 c net141 VSS VSS LPNFET W=0.44U L=0.12U M=1 
X39 VDD CK net141 VDD LPPFET W=0.34U L=0.12U M=1 
X4 hnet36 RN VSS VSS LPNFET W=0.98U L=0.12U M=1 
X40 net141 CK VSS VSS LPNFET W=0.34U L=0.12U M=1 
X5 m pm hnet36 VSS LPNFET W=0.98U L=0.12U M=1 
X6 net80 CK VDD VDD LPPFET W=0.98U L=0.12U M=1 
X7 cn c net80 VDD LPPFET W=0.74U L=0.12U M=1 
X8 nmsi SE nmin VDD LPPFET W=0.7U L=0.12U M=1 
X9 net122 RN VDD VDD LPPFET W=0.4U L=0.12U M=1 
.ENDS SDFFRHQX2TS 

**** 
*.SUBCKT SDFFRHQX4TS Q CK D RN SE SI 
.SUBCKT SDFFRHQX4TS Q CK D RN SE SI VSS VDD
X0 hnet29 cn VSS VSS LPNFET W=0.82U L=0.12U M=1 
X1 pm nmsi hnet29 VSS LPNFET W=0.82U L=0.12U M=1 
X10 VDD c hnet40 VDD LPPFET W=0.96U L=0.12U M=1 
X11 hnet40 nmsi pm VDD LPPFET W=0.96U L=0.12U M=1 
X12 net83 CK VDD VDD LPPFET W=0.84U L=0.12U M=1 
X13 cn c net83 VDD LPPFET W=0.64U L=0.12U M=1 
X14 net89 CK VDD VDD LPPFET W=0.84U L=0.12U M=1 
X15 cn c net89 VDD LPPFET W=0.64U L=0.12U M=1 
X16 nmsi SE nmin VDD LPPFET W=1.3U L=0.12U M=1 
X17 net131 RN VDD VDD LPPFET W=0.7U L=0.12U M=1 
X18 net131 c net100 VDD LPPFET W=0.28U L=0.12U M=1 
X19 net100 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X2 hnet33 cn VSS VSS LPNFET W=0.58U L=0.12U M=1 
X20 m RN VDD VDD LPPFET W=0.76U L=0.12U M=1 
X21 m pm VDD VDD LPPFET W=2.54U L=0.12U M=1 
X22 net131 cn m VDD LPPFET W=2.64U L=0.12U M=1 
X23 cn CK VSS VSS LPNFET W=0.48U L=0.12U M=1 
X24 nmsi nmse nmin VSS LPNFET W=0.84U L=0.12U M=1 
X25 net124 RN net121 VSS LPNFET W=0.2U L=0.12U M=1 
X26 net131 cn net124 VSS LPNFET W=0.2U L=0.12U M=1 
X27 net121 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X28 net131 c m VSS LPNFET W=1.4U L=0.12U M=1 
X29 hnet45 SI VSS VSS LPNFET W=0.46U L=0.12U M=1 
X3 pm nmsi hnet33 VSS LPNFET W=0.58U L=0.12U M=1 
X30 nmsi SE hnet45 VSS LPNFET W=0.46U L=0.12U M=1 
X31 hnet47 nmse nmsi VDD LPPFET W=0.66U L=0.12U M=1 
X32 VDD SI hnet47 VDD LPPFET W=0.66U L=0.12U M=1 
X33 hnet51 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X34 pm c hnet51 VSS LPNFET W=0.2U L=0.12U M=1 
X35 hnet53 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X36 VDD m hnet53 VDD LPPFET W=0.28U L=0.12U M=1 
X37 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X38 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X39 VDD D nmin VDD LPPFET W=1.3U L=0.12U M=1 
X4 hnet38 RN VSS VSS LPNFET W=0.8U L=0.12U M=1 
X40 nmin D VSS VSS LPNFET W=0.84U L=0.12U M=1 
X41 VDD net131 s VDD LPPFET W=0.28U L=0.12U M=1 
X42 s net131 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X43 VDD net131 Q VDD LPPFET W=2.6U L=0.12U M=1 
X44 Q net131 VSS VSS LPNFET W=1.66U L=0.12U M=1 
X45 VDD net150 c VDD LPPFET W=1.96U L=0.12U M=1 
X46 c net150 VSS VSS LPNFET W=0.72U L=0.12U M=1 
X47 VDD CK net150 VDD LPPFET W=0.56U L=0.12U M=1 
X48 net150 CK VSS VSS LPNFET W=0.56U L=0.12U M=1 
X5 m pm hnet38 VSS LPNFET W=0.8U L=0.12U M=1 
X6 hnet34 RN VSS VSS LPNFET W=0.8U L=0.12U M=1 
X7 m pm hnet34 VSS LPNFET W=0.8U L=0.12U M=1 
X8 VDD c hnet43 VDD LPPFET W=0.96U L=0.12U M=1 
X9 hnet43 nmsi pm VDD LPPFET W=0.96U L=0.12U M=1 
.ENDS SDFFRHQX4TS 

**** 
*.SUBCKT SDFFRHQX8TS Q CK D RN SE SI 
.SUBCKT SDFFRHQX8TS Q CK D RN SE SI VSS VDD
X0 hnet29 cn VSS VSS LPNFET W=0.82U L=0.12U M=1 
X1 pm nmsi hnet29 VSS LPNFET W=0.82U L=0.12U M=1 
X10 VDD c hnet40 VDD LPPFET W=0.96U L=0.12U M=1 
X11 hnet40 nmsi pm VDD LPPFET W=0.96U L=0.12U M=1 
X12 net85 CK VDD VDD LPPFET W=0.84U L=0.12U M=1 
X13 cn c net85 VDD LPPFET W=0.64U L=0.12U M=1 
X14 net91 CK VDD VDD LPPFET W=0.84U L=0.12U M=1 
X15 cn c net91 VDD LPPFET W=0.64U L=0.12U M=1 
X16 nmsi SE nmin VDD LPPFET W=1.3U L=0.12U M=1 
X17 net131 RN VDD VDD LPPFET W=0.7U L=0.12U M=1 
X18 net131 c net100 VDD LPPFET W=0.28U L=0.12U M=1 
X19 net100 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X2 hnet33 cn VSS VSS LPNFET W=0.58U L=0.12U M=1 
X20 m RN VDD VDD LPPFET W=0.76U L=0.12U M=1 
X21 m pm VDD VDD LPPFET W=2.54U L=0.12U M=1 
X22 net131 cn m VDD LPPFET W=2.64U L=0.12U M=1 
X23 cn CK VSS VSS LPNFET W=0.48U L=0.12U M=1 
X24 nmsi nmse nmin VSS LPNFET W=0.84U L=0.12U M=1 
X25 net124 RN net128 VSS LPNFET W=0.2U L=0.12U M=1 
X26 net131 cn net124 VSS LPNFET W=0.2U L=0.12U M=1 
X27 net128 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X28 net131 c m VSS LPNFET W=1.4U L=0.12U M=1 
X29 hnet45 SI VSS VSS LPNFET W=0.46U L=0.12U M=1 
X3 pm nmsi hnet33 VSS LPNFET W=0.58U L=0.12U M=1 
X30 nmsi SE hnet45 VSS LPNFET W=0.46U L=0.12U M=1 
X31 hnet47 nmse nmsi VDD LPPFET W=0.66U L=0.12U M=1 
X32 VDD SI hnet47 VDD LPPFET W=0.66U L=0.12U M=1 
X33 hnet51 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X34 pm c hnet51 VSS LPNFET W=0.2U L=0.12U M=1 
X35 hnet53 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X36 VDD m hnet53 VDD LPPFET W=0.28U L=0.12U M=1 
X37 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X38 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X39 VDD D nmin VDD LPPFET W=1.3U L=0.12U M=1 
X4 hnet38 RN VSS VSS LPNFET W=0.8U L=0.12U M=1 
X40 nmin D VSS VSS LPNFET W=0.84U L=0.12U M=1 
X41 VDD net131 s VDD LPPFET W=0.28U L=0.12U M=1 
X42 s net131 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X43 VDD net131 Q VDD LPPFET W=5.2U L=0.12U M=1 
X44 Q net131 VSS VSS LPNFET W=3.32U L=0.12U M=1 
X45 VDD net150 c VDD LPPFET W=1.96U L=0.12U M=1 
X46 c net150 VSS VSS LPNFET W=0.72U L=0.12U M=1 
X47 VDD CK net150 VDD LPPFET W=0.56U L=0.12U M=1 
X48 net150 CK VSS VSS LPNFET W=0.56U L=0.12U M=1 
X5 m pm hnet38 VSS LPNFET W=0.8U L=0.12U M=1 
X6 hnet34 RN VSS VSS LPNFET W=0.8U L=0.12U M=1 
X7 m pm hnet34 VSS LPNFET W=0.8U L=0.12U M=1 
X8 VDD c hnet43 VDD LPPFET W=0.96U L=0.12U M=1 
X9 hnet43 nmsi pm VDD LPPFET W=0.96U L=0.12U M=1 
.ENDS SDFFRHQX8TS 

**** 
*.SUBCKT SDFFRX1TS Q QN CK D RN SE SI 
.SUBCKT SDFFRX1TS Q QN CK D RN SE SI VSS VDD
X0 VDD D hnet29 VDD LPPFET W=0.36U L=0.12U M=1 
X1 hnet29 SE nmrs VDD LPPFET W=0.36U L=0.12U M=1 
X10 s net127 hnet47 VSS LPNFET W=0.32U L=0.12U M=1 
X11 VDD RN s VDD LPPFET W=0.28U L=0.12U M=1 
X12 VDD net127 s VDD LPPFET W=0.28U L=0.12U M=1 
X13 pm c nmrs VDD LPPFET W=0.28U L=0.12U M=1 
X14 pm RN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X15 net127 c net93 VDD LPPFET W=0.28U L=0.12U M=1 
X16 net93 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X17 net127 cn m VDD LPPFET W=0.28U L=0.12U M=1 
X18 net103 RN VSS VSS LPNFET W=0.44U L=0.12U M=1 
X19 net108 D net103 VSS LPNFET W=0.26U L=0.12U M=1 
X2 VDD SI hnet33 VDD LPPFET W=0.28U L=0.12U M=1 
X20 nmrs nmse net108 VSS LPNFET W=0.26U L=0.12U M=1 
X21 net114 SI net103 VSS LPNFET W=0.2U L=0.12U M=1 
X22 nmrs SE net114 VSS LPNFET W=0.2U L=0.12U M=1 
X23 pm cn nmrs VSS LPNFET W=0.2U L=0.12U M=1 
X24 net127 cn net124 VSS LPNFET W=0.2U L=0.12U M=1 
X25 net124 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X26 net127 c m VSS LPNFET W=0.2U L=0.12U M=1 
X27 VDD s net128 VDD LPPFET W=0.28U L=0.12U M=1 
X28 net128 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X29 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X3 hnet33 nmse nmrs VDD LPPFET W=0.28U L=0.12U M=1 
X30 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X31 VDD pm m VDD LPPFET W=0.28U L=0.12U M=1 
X32 m pm VSS VSS LPNFET W=0.2U L=0.12U M=1 
X33 VDD s Q VDD LPPFET W=0.64U L=0.12U M=1 
X34 Q s VSS VSS LPNFET W=0.46U L=0.12U M=1 
X35 VDD net128 QN VDD LPPFET W=0.64U L=0.12U M=1 
X36 QN net128 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X37 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X38 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X39 VDD CK cn VDD LPPFET W=0.42U L=0.12U M=1 
X4 VDD m hnet37 VDD LPPFET W=0.28U L=0.12U M=1 
X40 cn CK VSS VSS LPNFET W=0.3U L=0.12U M=1 
X5 hnet37 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X6 hnet43 RN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X7 hnet38 m hnet43 VSS LPNFET W=0.2U L=0.12U M=1 
X8 pm c hnet38 VSS LPNFET W=0.2U L=0.12U M=1 
X9 hnet47 RN VSS VSS LPNFET W=0.32U L=0.12U M=1 
.ENDS SDFFRX1TS 

**** 
*.SUBCKT SDFFRX2TS Q QN CK D RN SE SI 
.SUBCKT SDFFRX2TS Q QN CK D RN SE SI VSS VDD
X0 VDD D hnet29 VDD LPPFET W=0.36U L=0.12U M=1 
X1 hnet29 SE nmrs VDD LPPFET W=0.36U L=0.12U M=1 
X10 s net127 hnet47 VSS LPNFET W=0.52U L=0.12U M=1 
X11 VDD RN s VDD LPPFET W=0.38U L=0.12U M=1 
X12 VDD net127 s VDD LPPFET W=0.38U L=0.12U M=1 
X13 pm c nmrs VDD LPPFET W=0.28U L=0.12U M=1 
X14 pm RN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X15 net127 c net93 VDD LPPFET W=0.28U L=0.12U M=1 
X16 net93 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X17 net127 cn m VDD LPPFET W=0.28U L=0.12U M=1 
X18 net103 RN VSS VSS LPNFET W=0.44U L=0.12U M=1 
X19 net108 D net103 VSS LPNFET W=0.26U L=0.12U M=1 
X2 VDD SI hnet33 VDD LPPFET W=0.28U L=0.12U M=1 
X20 nmrs nmse net108 VSS LPNFET W=0.26U L=0.12U M=1 
X21 net112 SI net103 VSS LPNFET W=0.2U L=0.12U M=1 
X22 nmrs SE net112 VSS LPNFET W=0.2U L=0.12U M=1 
X23 pm cn nmrs VSS LPNFET W=0.2U L=0.12U M=1 
X24 net127 cn net124 VSS LPNFET W=0.2U L=0.12U M=1 
X25 net124 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X26 net127 c m VSS LPNFET W=0.2U L=0.12U M=1 
X27 VDD s net128 VDD LPPFET W=0.3U L=0.12U M=1 
X28 net128 s VSS VSS LPNFET W=0.22U L=0.12U M=1 
X29 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X3 hnet33 nmse nmrs VDD LPPFET W=0.28U L=0.12U M=1 
X30 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X31 VDD pm m VDD LPPFET W=0.28U L=0.12U M=1 
X32 m pm VSS VSS LPNFET W=0.2U L=0.12U M=1 
X33 VDD s Q VDD LPPFET W=1.28U L=0.12U M=1 
X34 Q s VSS VSS LPNFET W=0.92U L=0.12U M=1 
X35 VDD net128 QN VDD LPPFET W=1.28U L=0.12U M=1 
X36 QN net128 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X37 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X38 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X39 VDD CK cn VDD LPPFET W=0.42U L=0.12U M=1 
X4 VDD m hnet37 VDD LPPFET W=0.28U L=0.12U M=1 
X40 cn CK VSS VSS LPNFET W=0.3U L=0.12U M=1 
X5 hnet37 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X6 hnet43 RN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X7 hnet38 m hnet43 VSS LPNFET W=0.2U L=0.12U M=1 
X8 pm c hnet38 VSS LPNFET W=0.2U L=0.12U M=1 
X9 hnet47 RN VSS VSS LPNFET W=0.52U L=0.12U M=1 
.ENDS SDFFRX2TS 

**** 
*.SUBCKT SDFFRX4TS Q QN CK D RN SE SI 
.SUBCKT SDFFRX4TS Q QN CK D RN SE SI VSS VDD
X0 VDD D hnet29 VDD LPPFET W=0.36U L=0.12U M=1 
X1 hnet29 SE nmrs VDD LPPFET W=0.36U L=0.12U M=1 
X10 s net127 hnet47 VSS LPNFET W=0.92U L=0.12U M=1 
X11 VDD RN s VDD LPPFET W=0.68U L=0.12U M=1 
X12 VDD net127 s VDD LPPFET W=0.68U L=0.12U M=1 
X13 pm c nmrs VDD LPPFET W=0.28U L=0.12U M=1 
X14 pm RN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X15 net127 c net93 VDD LPPFET W=0.28U L=0.12U M=1 
X16 net93 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X17 net127 cn m VDD LPPFET W=0.48U L=0.12U M=1 
X18 net103 RN VSS VSS LPNFET W=0.44U L=0.12U M=1 
X19 net108 D net103 VSS LPNFET W=0.26U L=0.12U M=1 
X2 VDD SI hnet33 VDD LPPFET W=0.28U L=0.12U M=1 
X20 nmrs nmse net108 VSS LPNFET W=0.26U L=0.12U M=1 
X21 net114 SI net103 VSS LPNFET W=0.2U L=0.12U M=1 
X22 nmrs SE net114 VSS LPNFET W=0.2U L=0.12U M=1 
X23 pm cn nmrs VSS LPNFET W=0.2U L=0.12U M=1 
X24 net127 cn net124 VSS LPNFET W=0.2U L=0.12U M=1 
X25 net124 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X26 net127 c m VSS LPNFET W=0.34U L=0.12U M=1 
X27 VDD s net128 VDD LPPFET W=0.62U L=0.12U M=1 
X28 net128 s VSS VSS LPNFET W=0.44U L=0.12U M=1 
X29 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X3 hnet33 nmse nmrs VDD LPPFET W=0.28U L=0.12U M=1 
X30 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X31 VDD pm m VDD LPPFET W=0.48U L=0.12U M=1 
X32 m pm VSS VSS LPNFET W=0.34U L=0.12U M=1 
X33 VDD s Q VDD LPPFET W=2.56U L=0.12U M=1 
X34 Q s VSS VSS LPNFET W=1.84U L=0.12U M=1 
X35 VDD net128 QN VDD LPPFET W=2.56U L=0.12U M=1 
X36 QN net128 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X37 VDD cn c VDD LPPFET W=0.34U L=0.12U M=1 
X38 c cn VSS VSS LPNFET W=0.24U L=0.12U M=1 
X39 VDD CK cn VDD LPPFET W=0.52U L=0.12U M=1 
X4 VDD m hnet37 VDD LPPFET W=0.28U L=0.12U M=1 
X40 cn CK VSS VSS LPNFET W=0.38U L=0.12U M=1 
X5 hnet37 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X6 hnet43 RN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X7 hnet38 m hnet43 VSS LPNFET W=0.2U L=0.12U M=1 
X8 pm c hnet38 VSS LPNFET W=0.2U L=0.12U M=1 
X9 hnet47 RN VSS VSS LPNFET W=0.92U L=0.12U M=1 
.ENDS SDFFRX4TS 

**** 
*.SUBCKT SDFFRXLTS Q QN CK D RN SE SI 
.SUBCKT SDFFRXLTS Q QN CK D RN SE SI VSS VDD
X0 VDD D hnet29 VDD LPPFET W=0.36U L=0.12U M=1 
X1 hnet29 SE nmrs VDD LPPFET W=0.36U L=0.12U M=1 
X10 s net127 hnet47 VSS LPNFET W=0.22U L=0.12U M=1 
X11 VDD RN s VDD LPPFET W=0.28U L=0.12U M=1 
X12 VDD net127 s VDD LPPFET W=0.28U L=0.12U M=1 
X13 pm c nmrs VDD LPPFET W=0.28U L=0.12U M=1 
X14 pm RN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X15 net127 c net93 VDD LPPFET W=0.28U L=0.12U M=1 
X16 net93 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X17 net127 cn m VDD LPPFET W=0.28U L=0.12U M=1 
X18 net103 RN VSS VSS LPNFET W=0.44U L=0.12U M=1 
X19 net108 D net103 VSS LPNFET W=0.26U L=0.12U M=1 
X2 VDD SI hnet33 VDD LPPFET W=0.28U L=0.12U M=1 
X20 nmrs nmse net108 VSS LPNFET W=0.26U L=0.12U M=1 
X21 net114 SI net103 VSS LPNFET W=0.2U L=0.12U M=1 
X22 nmrs SE net114 VSS LPNFET W=0.2U L=0.12U M=1 
X23 pm cn nmrs VSS LPNFET W=0.2U L=0.12U M=1 
X24 net127 cn net124 VSS LPNFET W=0.2U L=0.12U M=1 
X25 net124 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X26 net127 c m VSS LPNFET W=0.2U L=0.12U M=1 
X27 VDD s net128 VDD LPPFET W=0.28U L=0.12U M=1 
X28 net128 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X29 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X3 hnet33 nmse nmrs VDD LPPFET W=0.28U L=0.12U M=1 
X30 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X31 VDD pm m VDD LPPFET W=0.28U L=0.12U M=1 
X32 m pm VSS VSS LPNFET W=0.2U L=0.12U M=1 
X33 VDD s Q VDD LPPFET W=0.34U L=0.12U M=1 
X34 Q s VSS VSS LPNFET W=0.24U L=0.12U M=1 
X35 VDD net128 QN VDD LPPFET W=0.34U L=0.12U M=1 
X36 QN net128 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X37 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X38 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X39 VDD CK cn VDD LPPFET W=0.42U L=0.12U M=1 
X4 VDD m hnet37 VDD LPPFET W=0.28U L=0.12U M=1 
X40 cn CK VSS VSS LPNFET W=0.3U L=0.12U M=1 
X5 hnet37 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X6 hnet43 RN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X7 hnet38 m hnet43 VSS LPNFET W=0.2U L=0.12U M=1 
X8 pm c hnet38 VSS LPNFET W=0.2U L=0.12U M=1 
X9 hnet47 RN VSS VSS LPNFET W=0.22U L=0.12U M=1 
.ENDS SDFFRXLTS 

**** 
*.SUBCKT SDFFSHQX1TS Q CK D SE SI SN 
.SUBCKT SDFFSHQX1TS Q CK D SE SI SN VSS VDD
X0 VDD c hnet29 VDD LPPFET W=0.52U L=0.12U M=1 
X1 hnet29 nmsi pm VDD LPPFET W=0.52U L=0.12U M=1 
X10 net112 c net87 VDD LPPFET W=0.26U L=0.12U M=1 
X11 net91 s VDD VDD LPPFET W=0.26U L=0.12U M=1 
X12 net112 cn m VDD LPPFET W=0.96U L=0.12U M=1 
X13 cn CK VSS VSS LPNFET W=0.2U L=0.12U M=1 
X14 nmsi nmse nmin VSS LPNFET W=0.3U L=0.12U M=1 
X15 net112 cn net106 VSS LPNFET W=0.2U L=0.12U M=1 
X16 net106 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X17 net112 nmset VSS VSS LPNFET W=0.2U L=0.12U M=1 
X18 net112 c m VSS LPNFET W=0.48U L=0.12U M=1 
X19 hnet37 SI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 hnet35 SN VSS VSS LPNFET W=0.54U L=0.12U M=1 
X20 nmsi SE hnet37 VSS LPNFET W=0.2U L=0.12U M=1 
X21 hnet39 nmse nmsi VDD LPPFET W=0.28U L=0.12U M=1 
X22 VDD SI hnet39 VDD LPPFET W=0.28U L=0.12U M=1 
X23 hnet43 m VSS VSS LPNFET W=0.18U L=0.12U M=1 
X24 pm c hnet43 VSS LPNFET W=0.18U L=0.12U M=1 
X25 hnet45 cn pm VDD LPPFET W=0.24U L=0.12U M=1 
X26 VDD m hnet45 VDD LPPFET W=0.24U L=0.12U M=1 
X27 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X28 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X29 VDD pm m VDD LPPFET W=0.96U L=0.12U M=1 
X3 hnet30 cn hnet35 VSS LPNFET W=0.54U L=0.12U M=1 
X30 m pm VSS VSS LPNFET W=0.46U L=0.12U M=1 
X31 VDD SN nmset VDD LPPFET W=0.28U L=0.12U M=1 
X32 nmset SN VSS VSS LPNFET W=0.18U L=0.12U M=1 
X33 VDD D nmin VDD LPPFET W=0.42U L=0.12U M=1 
X34 nmin D VSS VSS LPNFET W=0.3U L=0.12U M=1 
X35 VDD net112 s VDD LPPFET W=0.26U L=0.12U M=1 
X36 s net112 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X37 VDD net112 Q VDD LPPFET W=0.74U L=0.12U M=1 
X38 Q net112 VSS VSS LPNFET W=0.38U L=0.12U M=1 
X39 VDD net135 c VDD LPPFET W=0.72U L=0.12U M=1 
X4 pm nmsi hnet30 VSS LPNFET W=0.54U L=0.12U M=1 
X40 c net135 VSS VSS LPNFET W=0.26U L=0.12U M=1 
X41 VDD CK net135 VDD LPPFET W=0.28U L=0.12U M=1 
X42 net135 CK VSS VSS LPNFET W=0.28U L=0.12U M=1 
X5 net75 CK VDD VDD LPPFET W=0.62U L=0.12U M=1 
X6 cn c net75 VDD LPPFET W=0.52U L=0.12U M=1 
X7 nmsi SE nmin VDD LPPFET W=0.42U L=0.12U M=1 
X8 pm SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X9 net87 nmset net91 VDD LPPFET W=0.26U L=0.12U M=1 
.ENDS SDFFSHQX1TS 

**** 
*.SUBCKT SDFFSHQX2TS Q CK D SE SI SN 
.SUBCKT SDFFSHQX2TS Q CK D SE SI SN VSS VDD
X0 VDD c hnet29 VDD LPPFET W=0.9U L=0.12U M=1 
X1 hnet29 nmsi pm VDD LPPFET W=0.9U L=0.12U M=1 
X10 net112 c net87 VDD LPPFET W=0.26U L=0.12U M=1 
X11 net91 s VDD VDD LPPFET W=0.26U L=0.12U M=1 
X12 net112 cn m VDD LPPFET W=1.64U L=0.12U M=1 
X13 cn CK VSS VSS LPNFET W=0.3U L=0.12U M=1 
X14 nmsi nmse nmin VSS LPNFET W=0.52U L=0.12U M=1 
X15 net112 cn net102 VSS LPNFET W=0.2U L=0.12U M=1 
X16 net102 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X17 net112 nmset VSS VSS LPNFET W=0.28U L=0.12U M=1 
X18 net112 c m VSS LPNFET W=0.82U L=0.12U M=1 
X19 hnet37 SI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 hnet35 SN VSS VSS LPNFET W=0.86U L=0.12U M=1 
X20 nmsi SE hnet37 VSS LPNFET W=0.2U L=0.12U M=1 
X21 hnet39 nmse nmsi VDD LPPFET W=0.28U L=0.12U M=1 
X22 VDD SI hnet39 VDD LPPFET W=0.28U L=0.12U M=1 
X23 hnet43 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X24 pm c hnet43 VSS LPNFET W=0.2U L=0.12U M=1 
X25 hnet45 cn pm VDD LPPFET W=0.26U L=0.12U M=1 
X26 VDD m hnet45 VDD LPPFET W=0.26U L=0.12U M=1 
X27 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X28 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X29 VDD pm m VDD LPPFET W=1.64U L=0.12U M=1 
X3 hnet30 cn hnet35 VSS LPNFET W=0.86U L=0.12U M=1 
X30 m pm VSS VSS LPNFET W=0.84U L=0.12U M=1 
X31 VDD SN nmset VDD LPPFET W=0.28U L=0.12U M=1 
X32 nmset SN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X33 VDD D nmin VDD LPPFET W=0.76U L=0.12U M=1 
X34 nmin D VSS VSS LPNFET W=0.54U L=0.12U M=1 
X35 VDD net112 s VDD LPPFET W=0.28U L=0.12U M=1 
X36 s net112 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X37 VDD net112 Q VDD LPPFET W=1.3U L=0.12U M=1 
X38 Q net112 VSS VSS LPNFET W=0.84U L=0.12U M=1 
X39 VDD net135 c VDD LPPFET W=1.06U L=0.12U M=1 
X4 pm nmsi hnet30 VSS LPNFET W=0.86U L=0.12U M=1 
X40 c net135 VSS VSS LPNFET W=0.42U L=0.12U M=1 
X41 VDD CK net135 VDD LPPFET W=0.32U L=0.12U M=1 
X42 net135 CK VSS VSS LPNFET W=0.32U L=0.12U M=1 
X5 net75 CK VDD VDD LPPFET W=1.06U L=0.12U M=1 
X6 cn c net75 VDD LPPFET W=0.78U L=0.12U M=1 
X7 nmsi SE nmin VDD LPPFET W=0.76U L=0.12U M=1 
X8 pm SN VDD VDD LPPFET W=0.34U L=0.12U M=1 
X9 net87 nmset net91 VDD LPPFET W=0.26U L=0.12U M=1 
.ENDS SDFFSHQX2TS 

**** 
*.SUBCKT SDFFSHQX4TS Q CK D SE SI SN 
.SUBCKT SDFFSHQX4TS Q CK D SE SI SN VSS VDD
X0 hnet32 SN VSS VSS LPNFET W=0.84U L=0.12U M=1 
X1 hnet26 cn hnet32 VSS LPNFET W=0.84U L=0.12U M=1 
X10 net75 CK VDD VDD LPPFET W=1.84U L=0.12U M=1 
X11 cn c net75 VDD LPPFET W=1.3U L=0.12U M=1 
X12 nmsi SE nmin VDD LPPFET W=1.3U L=0.12U M=1 
X13 pm SN VDD VDD LPPFET W=0.64U L=0.12U M=1 
X14 net87 nmset net91 VDD LPPFET W=0.28U L=0.12U M=1 
X15 net112 c net87 VDD LPPFET W=0.28U L=0.12U M=1 
X16 net91 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X17 net112 cn m VDD LPPFET W=2.32U L=0.12U M=1 
X18 cn CK VSS VSS LPNFET W=0.52U L=0.12U M=1 
X19 nmsi nmse nmin VSS LPNFET W=0.92U L=0.12U M=1 
X2 pm nmsi hnet26 VSS LPNFET W=0.84U L=0.12U M=1 
X20 net112 cn net102 VSS LPNFET W=0.2U L=0.12U M=1 
X21 net102 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X22 net112 nmset VSS VSS LPNFET W=0.52U L=0.12U M=1 
X23 net112 c m VSS LPNFET W=1.36U L=0.12U M=1 
X24 hnet40 SI VSS VSS LPNFET W=0.34U L=0.12U M=1 
X25 nmsi SE hnet40 VSS LPNFET W=0.34U L=0.12U M=1 
X26 hnet42 nmse nmsi VDD LPPFET W=0.48U L=0.12U M=1 
X27 VDD SI hnet42 VDD LPPFET W=0.48U L=0.12U M=1 
X28 hnet46 m VSS VSS LPNFET W=0.22U L=0.12U M=1 
X29 pm c hnet46 VSS LPNFET W=0.22U L=0.12U M=1 
X3 hnet33 SN VSS VSS LPNFET W=0.84U L=0.12U M=1 
X30 hnet48 cn pm VDD LPPFET W=0.3U L=0.12U M=1 
X31 VDD m hnet48 VDD LPPFET W=0.3U L=0.12U M=1 
X32 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X33 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X34 VDD pm m VDD LPPFET W=3U L=0.12U M=1 
X35 m pm VSS VSS LPNFET W=1.48U L=0.12U M=1 
X36 VDD SN nmset VDD LPPFET W=0.28U L=0.12U M=1 
X37 nmset SN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X38 VDD D nmin VDD LPPFET W=1.34U L=0.12U M=1 
X39 nmin D VSS VSS LPNFET W=0.92U L=0.12U M=1 
X4 hnet28 cn hnet33 VSS LPNFET W=0.84U L=0.12U M=1 
X40 VDD net112 s VDD LPPFET W=0.28U L=0.12U M=1 
X41 s net112 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X42 VDD net112 Q VDD LPPFET W=2.6U L=0.12U M=1 
X43 Q net112 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X44 VDD net135 c VDD LPPFET W=2.02U L=0.12U M=1 
X45 c net135 VSS VSS LPNFET W=0.72U L=0.12U M=1 
X46 VDD CK net135 VDD LPPFET W=0.54U L=0.12U M=1 
X47 net135 CK VSS VSS LPNFET W=0.54U L=0.12U M=1 
X5 pm nmsi hnet28 VSS LPNFET W=0.84U L=0.12U M=1 
X6 VDD c hnet38 VDD LPPFET W=0.74U L=0.12U M=1 
X7 hnet38 nmsi pm VDD LPPFET W=0.74U L=0.12U M=1 
X8 VDD c hnet35 VDD LPPFET W=0.74U L=0.12U M=1 
X9 hnet35 nmsi pm VDD LPPFET W=0.74U L=0.12U M=1 
.ENDS SDFFSHQX4TS 

**** 
*.SUBCKT SDFFSHQX8TS Q CK D SE SI SN 
.SUBCKT SDFFSHQX8TS Q CK D SE SI SN VSS VDD
X0 hnet32 SN VSS VSS LPNFET W=0.84U L=0.12U M=1 
X1 hnet26 cn hnet32 VSS LPNFET W=0.84U L=0.12U M=1 
X10 net75 CK VDD VDD LPPFET W=1.84U L=0.12U M=1 
X11 cn c net75 VDD LPPFET W=1.3U L=0.12U M=1 
X12 nmsi SE nmin VDD LPPFET W=1.3U L=0.12U M=1 
X13 pm SN VDD VDD LPPFET W=0.64U L=0.12U M=1 
X14 net87 nmset net91 VDD LPPFET W=0.28U L=0.12U M=1 
X15 net112 c net87 VDD LPPFET W=0.28U L=0.12U M=1 
X16 net91 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X17 net112 cn m VDD LPPFET W=2.3U L=0.12U M=1 
X18 cn CK VSS VSS LPNFET W=0.52U L=0.12U M=1 
X19 nmsi nmse nmin VSS LPNFET W=0.92U L=0.12U M=1 
X2 pm nmsi hnet26 VSS LPNFET W=0.84U L=0.12U M=1 
X20 net112 cn net102 VSS LPNFET W=0.2U L=0.12U M=1 
X21 net102 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X22 net112 nmset VSS VSS LPNFET W=0.52U L=0.12U M=1 
X23 net112 c m VSS LPNFET W=1.36U L=0.12U M=1 
X24 hnet40 SI VSS VSS LPNFET W=0.34U L=0.12U M=1 
X25 nmsi SE hnet40 VSS LPNFET W=0.34U L=0.12U M=1 
X26 hnet42 nmse nmsi VDD LPPFET W=0.48U L=0.12U M=1 
X27 VDD SI hnet42 VDD LPPFET W=0.48U L=0.12U M=1 
X28 hnet46 m VSS VSS LPNFET W=0.22U L=0.12U M=1 
X29 pm c hnet46 VSS LPNFET W=0.22U L=0.12U M=1 
X3 hnet33 SN VSS VSS LPNFET W=0.84U L=0.12U M=1 
X30 hnet48 cn pm VDD LPPFET W=0.3U L=0.12U M=1 
X31 VDD m hnet48 VDD LPPFET W=0.3U L=0.12U M=1 
X32 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X33 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X34 VDD pm m VDD LPPFET W=3.12U L=0.12U M=1 
X35 m pm VSS VSS LPNFET W=1.48U L=0.12U M=1 
X36 VDD SN nmset VDD LPPFET W=0.28U L=0.12U M=1 
X37 nmset SN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X38 VDD D nmin VDD LPPFET W=1.34U L=0.12U M=1 
X39 nmin D VSS VSS LPNFET W=0.92U L=0.12U M=1 
X4 hnet28 cn hnet33 VSS LPNFET W=0.84U L=0.12U M=1 
X40 VDD net112 s VDD LPPFET W=0.28U L=0.12U M=1 
X41 s net112 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X42 VDD net112 Q VDD LPPFET W=5.2U L=0.12U M=1 
X43 Q net112 VSS VSS LPNFET W=3.68U L=0.12U M=1 
X44 VDD net135 c VDD LPPFET W=2U L=0.12U M=1 
X45 c net135 VSS VSS LPNFET W=0.72U L=0.12U M=1 
X46 VDD CK net135 VDD LPPFET W=0.54U L=0.12U M=1 
X47 net135 CK VSS VSS LPNFET W=0.54U L=0.12U M=1 
X5 pm nmsi hnet28 VSS LPNFET W=0.84U L=0.12U M=1 
X6 VDD c hnet38 VDD LPPFET W=0.74U L=0.12U M=1 
X7 hnet38 nmsi pm VDD LPPFET W=0.74U L=0.12U M=1 
X8 VDD c hnet35 VDD LPPFET W=0.74U L=0.12U M=1 
X9 hnet35 nmsi pm VDD LPPFET W=0.74U L=0.12U M=1 
.ENDS SDFFSHQX8TS 

**** 
*.SUBCKT SDFFSRHQX1TS Q CK D RN SE SI SN 
.SUBCKT SDFFSRHQX1TS Q CK D RN SE SI SN VSS VDD
X0 hnet33 SN VSS VSS LPNFET W=0.54U L=0.12U M=1 
X1 hnet28 cn hnet33 VSS LPNFET W=0.54U L=0.12U M=1 
X10 hnet49 nmset net148 VDD LPPFET W=0.28U L=0.12U M=1 
X11 net102 CK VDD VDD LPPFET W=0.7U L=0.12U M=1 
X12 cn c net102 VDD LPPFET W=0.52U L=0.12U M=1 
X13 nmsi SE nmin VDD LPPFET W=0.38U L=0.12U M=1 
X14 pm SN VDD VDD LPPFET W=0.26U L=0.12U M=1 
X15 m pm VDD VDD LPPFET W=0.66U L=0.12U M=1 
X16 net115 nmset net121 VDD LPPFET W=0.26U L=0.12U M=1 
X17 net148 c net115 VDD LPPFET W=0.26U L=0.12U M=1 
X18 net121 s VDD VDD LPPFET W=0.26U L=0.12U M=1 
X19 net148 cn m VDD LPPFET W=0.66U L=0.12U M=1 
X2 pm nmsi hnet28 VSS LPNFET W=0.54U L=0.12U M=1 
X20 cn CK VSS VSS LPNFET W=0.2U L=0.12U M=1 
X21 nmsi nmse nmin VSS LPNFET W=0.28U L=0.12U M=1 
X22 net133 RN net132 VSS LPNFET W=0.2U L=0.12U M=1 
X23 net148 cn net133 VSS LPNFET W=0.2U L=0.12U M=1 
X24 net132 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X25 net148 nmset VSS VSS LPNFET W=0.2U L=0.12U M=1 
X26 m nmset VSS VSS LPNFET W=0.2U L=0.12U M=1 
X27 net148 c m VSS LPNFET W=0.46U L=0.12U M=1 
X28 hnet51 SI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X29 nmsi SE hnet51 VSS LPNFET W=0.2U L=0.12U M=1 
X3 hnet37 RN VSS VSS LPNFET W=0.5U L=0.12U M=1 
X30 hnet53 nmse nmsi VDD LPPFET W=0.28U L=0.12U M=1 
X31 VDD SI hnet53 VDD LPPFET W=0.28U L=0.12U M=1 
X32 hnet57 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X33 pm c hnet57 VSS LPNFET W=0.2U L=0.12U M=1 
X34 hnet59 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X35 VDD m hnet59 VDD LPPFET W=0.28U L=0.12U M=1 
X36 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X37 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X38 VDD SN nmset VDD LPPFET W=0.28U L=0.12U M=1 
X39 nmset SN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X4 m pm hnet37 VSS LPNFET W=0.5U L=0.12U M=1 
X40 VDD D nmin VDD LPPFET W=0.38U L=0.12U M=1 
X41 nmin D VSS VSS LPNFET W=0.28U L=0.12U M=1 
X42 VDD net148 s VDD LPPFET W=0.28U L=0.12U M=1 
X43 s net148 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X44 VDD net148 Q VDD LPPFET W=0.76U L=0.12U M=1 
X45 Q net148 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X46 VDD net169 c VDD LPPFET W=0.78U L=0.12U M=1 
X47 c net169 VSS VSS LPNFET W=0.28U L=0.12U M=1 
X48 VDD CK net169 VDD LPPFET W=0.28U L=0.12U M=1 
X49 net169 CK VSS VSS LPNFET W=0.28U L=0.12U M=1 
X5 VDD c hnet41 VDD LPPFET W=0.46U L=0.12U M=1 
X6 hnet41 nmsi pm VDD LPPFET W=0.46U L=0.12U M=1 
X7 VDD nmset hnet45 VDD LPPFET W=0.26U L=0.12U M=1 
X8 hnet45 RN m VDD LPPFET W=0.26U L=0.12U M=1 
X9 VDD RN hnet49 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS SDFFSRHQX1TS 

**** 
*.SUBCKT SDFFSRHQX2TS Q CK D RN SE SI SN 
.SUBCKT SDFFSRHQX2TS Q CK D RN SE SI SN VSS VDD
X0 hnet33 SN VSS VSS LPNFET W=0.88U L=0.12U M=1 
X1 hnet28 cn hnet33 VSS LPNFET W=0.88U L=0.12U M=1 
X10 hnet49 nmset net148 VDD LPPFET W=0.46U L=0.12U M=1 
X11 net102 CK VDD VDD LPPFET W=0.86U L=0.12U M=1 
X12 cn c net102 VDD LPPFET W=0.64U L=0.12U M=1 
X13 nmsi SE nmin VDD LPPFET W=0.7U L=0.12U M=1 
X14 pm SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X15 m pm VDD VDD LPPFET W=1.14U L=0.12U M=1 
X16 net117 nmset net121 VDD LPPFET W=0.28U L=0.12U M=1 
X17 net148 c net117 VDD LPPFET W=0.28U L=0.12U M=1 
X18 net121 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X19 net148 cn m VDD LPPFET W=1.14U L=0.12U M=1 
X2 pm nmsi hnet28 VSS LPNFET W=0.88U L=0.12U M=1 
X20 cn CK VSS VSS LPNFET W=0.24U L=0.12U M=1 
X21 nmsi nmse nmin VSS LPNFET W=0.5U L=0.12U M=1 
X22 net135 RN net139 VSS LPNFET W=0.2U L=0.12U M=1 
X23 net148 cn net135 VSS LPNFET W=0.2U L=0.12U M=1 
X24 net139 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X25 net148 nmset VSS VSS LPNFET W=0.2U L=0.12U M=1 
X26 m nmset VSS VSS LPNFET W=0.2U L=0.12U M=1 
X27 net148 c m VSS LPNFET W=0.82U L=0.12U M=1 
X28 hnet51 SI VSS VSS LPNFET W=0.24U L=0.12U M=1 
X29 nmsi SE hnet51 VSS LPNFET W=0.24U L=0.12U M=1 
X3 hnet37 RN VSS VSS LPNFET W=0.86U L=0.12U M=1 
X30 hnet53 nmse nmsi VDD LPPFET W=0.34U L=0.12U M=1 
X31 VDD SI hnet53 VDD LPPFET W=0.34U L=0.12U M=1 
X32 hnet57 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X33 pm c hnet57 VSS LPNFET W=0.2U L=0.12U M=1 
X34 hnet59 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X35 VDD m hnet59 VDD LPPFET W=0.28U L=0.12U M=1 
X36 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X37 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X38 VDD SN nmset VDD LPPFET W=0.28U L=0.12U M=1 
X39 nmset SN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X4 m pm hnet37 VSS LPNFET W=0.86U L=0.12U M=1 
X40 VDD D nmin VDD LPPFET W=0.7U L=0.12U M=1 
X41 nmin D VSS VSS LPNFET W=0.5U L=0.12U M=1 
X42 VDD net148 s VDD LPPFET W=0.28U L=0.12U M=1 
X43 s net148 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X44 VDD net148 Q VDD LPPFET W=1.48U L=0.12U M=1 
X45 Q net148 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X46 VDD net169 c VDD LPPFET W=1.1U L=0.12U M=1 
X47 c net169 VSS VSS LPNFET W=0.4U L=0.12U M=1 
X48 VDD CK net169 VDD LPPFET W=0.3U L=0.12U M=1 
X49 net169 CK VSS VSS LPNFET W=0.3U L=0.12U M=1 
X5 VDD c hnet41 VDD LPPFET W=0.8U L=0.12U M=1 
X6 hnet41 nmsi pm VDD LPPFET W=0.8U L=0.12U M=1 
X7 VDD nmset hnet45 VDD LPPFET W=0.28U L=0.12U M=1 
X8 hnet45 RN m VDD LPPFET W=0.28U L=0.12U M=1 
X9 VDD RN hnet49 VDD LPPFET W=0.46U L=0.12U M=1 
.ENDS SDFFSRHQX2TS 

**** 
*.SUBCKT SDFFSRHQX4TS Q CK D RN SE SI SN 
.SUBCKT SDFFSRHQX4TS Q CK D RN SE SI SN VSS VDD
X0 hnet34 SN VSS VSS LPNFET W=1.1U L=0.12U M=1 
X1 hnet29 cn hnet34 VSS LPNFET W=1.1U L=0.12U M=1 
X10 hnet41 nmsi pm VDD LPPFET W=0.68U L=0.12U M=1 
X11 VDD nmset hnet48 VDD LPPFET W=0.52U L=0.12U M=1 
X12 hnet48 RN m VDD LPPFET W=0.52U L=0.12U M=1 
X13 VDD RN hnet52 VDD LPPFET W=0.84U L=0.12U M=1 
X14 hnet52 nmset net156 VDD LPPFET W=0.84U L=0.12U M=1 
X15 net110 CK VDD VDD LPPFET W=0.74U L=0.12U M=1 
X16 cn c net104 VDD LPPFET W=0.56U L=0.12U M=1 
X17 net104 CK VDD VDD LPPFET W=0.74U L=0.12U M=1 
X18 cn c net110 VDD LPPFET W=0.56U L=0.12U M=1 
X19 nmsi SE nmin VDD LPPFET W=1.24U L=0.12U M=1 
X2 pm nmsi hnet29 VSS LPNFET W=1.1U L=0.12U M=1 
X20 pm SN VDD VDD LPPFET W=0.36U L=0.12U M=1 
X21 m pm VDD VDD LPPFET W=2.08U L=0.12U M=1 
X22 net125 nmset net129 VDD LPPFET W=0.28U L=0.12U M=1 
X23 net156 c net125 VDD LPPFET W=0.28U L=0.12U M=1 
X24 net129 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X25 net156 cn m VDD LPPFET W=1.28U L=0.12U M=1 
X26 cn CK VSS VSS LPNFET W=0.42U L=0.12U M=1 
X27 nmsi nmse nmin VSS LPNFET W=0.86U L=0.12U M=1 
X28 net143 RN net147 VSS LPNFET W=0.2U L=0.12U M=1 
X29 net156 cn net143 VSS LPNFET W=0.2U L=0.12U M=1 
X3 hnet39 RN VSS VSS LPNFET W=0.5U L=0.12U M=1 
X30 net147 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X31 net156 nmset VSS VSS LPNFET W=0.38U L=0.12U M=1 
X32 m nmset VSS VSS LPNFET W=0.38U L=0.12U M=1 
X33 net156 c m VSS LPNFET W=0.92U L=0.12U M=1 
X34 hnet54 SI VSS VSS LPNFET W=0.44U L=0.12U M=1 
X35 nmsi SE hnet54 VSS LPNFET W=0.44U L=0.12U M=1 
X36 hnet56 nmse nmsi VDD LPPFET W=0.62U L=0.12U M=1 
X37 VDD SI hnet56 VDD LPPFET W=0.62U L=0.12U M=1 
X38 hnet60 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X39 pm c hnet60 VSS LPNFET W=0.2U L=0.12U M=1 
X4 m pm hnet39 VSS LPNFET W=0.5U L=0.12U M=1 
X40 hnet62 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X41 VDD m hnet62 VDD LPPFET W=0.28U L=0.12U M=1 
X42 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X43 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X44 VDD SN nmset VDD LPPFET W=0.34U L=0.12U M=1 
X45 nmset SN VSS VSS LPNFET W=0.24U L=0.12U M=1 
X46 VDD D nmin VDD LPPFET W=1.24U L=0.12U M=1 
X47 nmin D VSS VSS LPNFET W=0.86U L=0.12U M=1 
X48 VDD net156 s VDD LPPFET W=0.28U L=0.12U M=1 
X49 s net156 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X5 hnet35 RN VSS VSS LPNFET W=0.5U L=0.12U M=1 
X50 VDD net156 Q VDD LPPFET W=2.6U L=0.12U M=1 
X51 Q net156 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X52 VDD net177 c VDD LPPFET W=1.66U L=0.12U M=1 
X53 c net177 VSS VSS LPNFET W=0.66U L=0.12U M=1 
X54 VDD CK net177 VDD LPPFET W=0.5U L=0.12U M=1 
X55 net177 CK VSS VSS LPNFET W=0.5U L=0.12U M=1 
X6 m pm hnet35 VSS LPNFET W=0.5U L=0.12U M=1 
X7 VDD c hnet44 VDD LPPFET W=0.68U L=0.12U M=1 
X8 hnet44 nmsi pm VDD LPPFET W=0.68U L=0.12U M=1 
X9 VDD c hnet41 VDD LPPFET W=0.68U L=0.12U M=1 
.ENDS SDFFSRHQX4TS 

**** 
*.SUBCKT SDFFSRHQX8TS Q CK D RN SE SI SN 
.SUBCKT SDFFSRHQX8TS Q CK D RN SE SI SN VSS VDD
X0 hnet34 SN VSS VSS LPNFET W=1.1U L=0.12U M=1 
X1 hnet29 cn hnet34 VSS LPNFET W=1.1U L=0.12U M=1 
X10 hnet41 nmsi pm VDD LPPFET W=0.68U L=0.12U M=1 
X11 VDD nmset hnet48 VDD LPPFET W=0.52U L=0.12U M=1 
X12 hnet48 RN m VDD LPPFET W=0.52U L=0.12U M=1 
X13 VDD RN hnet52 VDD LPPFET W=0.84U L=0.12U M=1 
X14 hnet52 nmset net156 VDD LPPFET W=0.84U L=0.12U M=1 
X15 net110 CK VDD VDD LPPFET W=0.74U L=0.12U M=1 
X16 cn c net104 VDD LPPFET W=0.56U L=0.12U M=1 
X17 net104 CK VDD VDD LPPFET W=0.74U L=0.12U M=1 
X18 cn c net110 VDD LPPFET W=0.56U L=0.12U M=1 
X19 nmsi SE nmin VDD LPPFET W=1.24U L=0.12U M=1 
X2 pm nmsi hnet29 VSS LPNFET W=1.1U L=0.12U M=1 
X20 pm SN VDD VDD LPPFET W=0.36U L=0.12U M=1 
X21 m pm VDD VDD LPPFET W=2.08U L=0.12U M=1 
X22 net125 nmset net129 VDD LPPFET W=0.28U L=0.12U M=1 
X23 net156 c net125 VDD LPPFET W=0.28U L=0.12U M=1 
X24 net129 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X25 net156 cn m VDD LPPFET W=1.28U L=0.12U M=1 
X26 cn CK VSS VSS LPNFET W=0.42U L=0.12U M=1 
X27 nmsi nmse nmin VSS LPNFET W=0.86U L=0.12U M=1 
X28 net143 RN net147 VSS LPNFET W=0.2U L=0.12U M=1 
X29 net156 cn net143 VSS LPNFET W=0.2U L=0.12U M=1 
X3 hnet39 RN VSS VSS LPNFET W=0.5U L=0.12U M=1 
X30 net147 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X31 net156 nmset VSS VSS LPNFET W=0.38U L=0.12U M=1 
X32 m nmset VSS VSS LPNFET W=0.38U L=0.12U M=1 
X33 net156 c m VSS LPNFET W=0.92U L=0.12U M=1 
X34 hnet54 SI VSS VSS LPNFET W=0.44U L=0.12U M=1 
X35 nmsi SE hnet54 VSS LPNFET W=0.44U L=0.12U M=1 
X36 hnet56 nmse nmsi VDD LPPFET W=0.62U L=0.12U M=1 
X37 VDD SI hnet56 VDD LPPFET W=0.62U L=0.12U M=1 
X38 hnet60 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X39 pm c hnet60 VSS LPNFET W=0.2U L=0.12U M=1 
X4 m pm hnet39 VSS LPNFET W=0.5U L=0.12U M=1 
X40 hnet62 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X41 VDD m hnet62 VDD LPPFET W=0.28U L=0.12U M=1 
X42 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X43 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X44 VDD SN nmset VDD LPPFET W=0.34U L=0.12U M=1 
X45 nmset SN VSS VSS LPNFET W=0.24U L=0.12U M=1 
X46 VDD D nmin VDD LPPFET W=1.24U L=0.12U M=1 
X47 nmin D VSS VSS LPNFET W=0.86U L=0.12U M=1 
X48 VDD net156 s VDD LPPFET W=0.28U L=0.12U M=1 
X49 s net156 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X5 hnet35 RN VSS VSS LPNFET W=0.5U L=0.12U M=1 
X50 VDD net156 Q VDD LPPFET W=5.2U L=0.12U M=1 
X51 Q net156 VSS VSS LPNFET W=3.68U L=0.12U M=1 
X52 VDD net177 c VDD LPPFET W=1.66U L=0.12U M=1 
X53 c net177 VSS VSS LPNFET W=0.66U L=0.12U M=1 
X54 VDD CK net177 VDD LPPFET W=0.5U L=0.12U M=1 
X55 net177 CK VSS VSS LPNFET W=0.5U L=0.12U M=1 
X6 m pm hnet35 VSS LPNFET W=0.5U L=0.12U M=1 
X7 VDD c hnet44 VDD LPPFET W=0.68U L=0.12U M=1 
X8 hnet44 nmsi pm VDD LPPFET W=0.68U L=0.12U M=1 
X9 VDD c hnet41 VDD LPPFET W=0.68U L=0.12U M=1 
.ENDS SDFFSRHQX8TS 

**** 
*.SUBCKT SDFFSRX1TS Q QN CK D RN SE SI SN 
.SUBCKT SDFFSRX1TS Q QN CK D RN SE SI SN VSS VDD
X0 VDD D hnet32 VDD LPPFET W=0.28U L=0.12U M=1 
X1 hnet32 SE nminsi VDD LPPFET W=0.28U L=0.12U M=1 
X10 net146 c net104 VDD LPPFET W=0.28U L=0.12U M=1 
X11 net146 cn m VDD LPPFET W=0.28U L=0.12U M=1 
X12 net115 D VSS VSS LPNFET W=0.2U L=0.12U M=1 
X13 nminsi nmse net115 VSS LPNFET W=0.2U L=0.12U M=1 
X14 net119 SI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X15 nminsi SE net119 VSS LPNFET W=0.2U L=0.12U M=1 
X16 pm cn nminsi VSS LPNFET W=0.2U L=0.12U M=1 
X17 m net157 net140 VSS LPNFET W=0.2U L=0.12U M=1 
X18 m pm net140 VSS LPNFET W=0.3U L=0.12U M=1 
X19 net146 net157 net140 VSS LPNFET W=0.2U L=0.12U M=1 
X2 VDD SI hnet36 VDD LPPFET W=0.28U L=0.12U M=1 
X20 net137 s net140 VSS LPNFET W=0.2U L=0.12U M=1 
X21 net140 SN VSS VSS LPNFET W=0.4U L=0.12U M=1 
X22 net146 cn net137 VSS LPNFET W=0.2U L=0.12U M=1 
X23 net146 c m VSS LPNFET W=0.2U L=0.12U M=1 
X24 hnet38 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X25 pm c hnet38 VSS LPNFET W=0.2U L=0.12U M=1 
X26 hnet40 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X27 VDD m hnet40 VDD LPPFET W=0.28U L=0.12U M=1 
X28 VDD s net151 VDD LPPFET W=0.28U L=0.12U M=1 
X29 net151 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 hnet36 nmse nminsi VDD LPPFET W=0.28U L=0.12U M=1 
X30 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X31 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X32 VDD s Q VDD LPPFET W=0.64U L=0.12U M=1 
X33 Q s VSS VSS LPNFET W=0.46U L=0.12U M=1 
X34 VDD RN net157 VDD LPPFET W=0.28U L=0.12U M=1 
X35 net157 RN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X36 VDD net146 s VDD LPPFET W=0.28U L=0.12U M=1 
X37 s net146 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X38 VDD net151 QN VDD LPPFET W=0.64U L=0.12U M=1 
X39 QN net151 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X4 pm c nminsi VDD LPPFET W=0.28U L=0.12U M=1 
X40 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X41 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X42 VDD CK cn VDD LPPFET W=0.42U L=0.12U M=1 
X43 cn CK VSS VSS LPNFET W=0.3U L=0.12U M=1 
X5 m SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X6 m pm net94 VDD LPPFET W=0.42U L=0.12U M=1 
X7 net94 net157 VDD VDD LPPFET W=0.56U L=0.12U M=1 
X8 net146 SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X9 net104 s net94 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS SDFFSRX1TS 

**** 
*.SUBCKT SDFFSRX2TS Q QN CK D RN SE SI SN 
.SUBCKT SDFFSRX2TS Q QN CK D RN SE SI SN VSS VDD
X0 VDD D hnet32 VDD LPPFET W=0.28U L=0.12U M=1 
X1 hnet32 SE nminsi VDD LPPFET W=0.28U L=0.12U M=1 
X10 net146 c net104 VDD LPPFET W=0.28U L=0.12U M=1 
X11 net146 cn m VDD LPPFET W=0.28U L=0.12U M=1 
X12 net115 D VSS VSS LPNFET W=0.2U L=0.12U M=1 
X13 nminsi nmse net115 VSS LPNFET W=0.2U L=0.12U M=1 
X14 net121 SI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X15 nminsi SE net121 VSS LPNFET W=0.2U L=0.12U M=1 
X16 pm cn nminsi VSS LPNFET W=0.2U L=0.12U M=1 
X17 m net157 net140 VSS LPNFET W=0.2U L=0.12U M=1 
X18 m pm net140 VSS LPNFET W=0.3U L=0.12U M=1 
X19 net146 net157 net140 VSS LPNFET W=0.2U L=0.12U M=1 
X2 VDD SI hnet36 VDD LPPFET W=0.28U L=0.12U M=1 
X20 net142 s net140 VSS LPNFET W=0.2U L=0.12U M=1 
X21 net140 SN VSS VSS LPNFET W=0.4U L=0.12U M=1 
X22 net146 cn net142 VSS LPNFET W=0.2U L=0.12U M=1 
X23 net146 c m VSS LPNFET W=0.2U L=0.12U M=1 
X24 hnet38 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X25 pm c hnet38 VSS LPNFET W=0.2U L=0.12U M=1 
X26 hnet40 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X27 VDD m hnet40 VDD LPPFET W=0.28U L=0.12U M=1 
X28 VDD s net151 VDD LPPFET W=0.3U L=0.12U M=1 
X29 net151 s VSS VSS LPNFET W=0.22U L=0.12U M=1 
X3 hnet36 nmse nminsi VDD LPPFET W=0.28U L=0.12U M=1 
X30 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X31 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X32 VDD s Q VDD LPPFET W=1.28U L=0.12U M=1 
X33 Q s VSS VSS LPNFET W=0.92U L=0.12U M=1 
X34 VDD RN net157 VDD LPPFET W=0.28U L=0.12U M=1 
X35 net157 RN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X36 VDD net146 s VDD LPPFET W=0.34U L=0.12U M=1 
X37 s net146 VSS VSS LPNFET W=0.28U L=0.12U M=1 
X38 VDD net151 QN VDD LPPFET W=1.28U L=0.12U M=1 
X39 QN net151 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X4 pm c nminsi VDD LPPFET W=0.28U L=0.12U M=1 
X40 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X41 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X42 VDD CK cn VDD LPPFET W=0.42U L=0.12U M=1 
X43 cn CK VSS VSS LPNFET W=0.3U L=0.12U M=1 
X5 m SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X6 m pm net94 VDD LPPFET W=0.42U L=0.12U M=1 
X7 net94 net157 VDD VDD LPPFET W=0.56U L=0.12U M=1 
X8 net146 SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X9 net104 s net94 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS SDFFSRX2TS 

**** 
*.SUBCKT SDFFSRX4TS Q QN CK D RN SE SI SN 
.SUBCKT SDFFSRX4TS Q QN CK D RN SE SI SN VSS VDD
X0 VDD D hnet32 VDD LPPFET W=0.28U L=0.12U M=1 
X1 hnet32 SE nminsi VDD LPPFET W=0.28U L=0.12U M=1 
X10 net146 c net104 VDD LPPFET W=0.28U L=0.12U M=1 
X11 net146 cn m VDD LPPFET W=0.3U L=0.12U M=1 
X12 net115 D VSS VSS LPNFET W=0.2U L=0.12U M=1 
X13 nminsi nmse net115 VSS LPNFET W=0.2U L=0.12U M=1 
X14 net121 SI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X15 nminsi SE net121 VSS LPNFET W=0.2U L=0.12U M=1 
X16 pm cn nminsi VSS LPNFET W=0.2U L=0.12U M=1 
X17 m net157 net140 VSS LPNFET W=0.2U L=0.12U M=1 
X18 m pm net140 VSS LPNFET W=0.34U L=0.12U M=1 
X19 net146 net157 net140 VSS LPNFET W=0.2U L=0.12U M=1 
X2 VDD SI hnet36 VDD LPPFET W=0.28U L=0.12U M=1 
X20 net142 s net140 VSS LPNFET W=0.2U L=0.12U M=1 
X21 net140 SN VSS VSS LPNFET W=0.46U L=0.12U M=1 
X22 net146 cn net142 VSS LPNFET W=0.2U L=0.12U M=1 
X23 net146 c m VSS LPNFET W=0.22U L=0.12U M=1 
X24 hnet38 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X25 pm c hnet38 VSS LPNFET W=0.2U L=0.12U M=1 
X26 hnet40 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X27 VDD m hnet40 VDD LPPFET W=0.28U L=0.12U M=1 
X28 VDD s net151 VDD LPPFET W=0.62U L=0.12U M=1 
X29 net151 s VSS VSS LPNFET W=0.4U L=0.12U M=1 
X3 hnet36 nmse nminsi VDD LPPFET W=0.28U L=0.12U M=1 
X30 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X31 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X32 VDD s Q VDD LPPFET W=2.4U L=0.12U M=1 
X33 Q s VSS VSS LPNFET W=1.84U L=0.12U M=1 
X34 VDD RN net157 VDD LPPFET W=0.28U L=0.12U M=1 
X35 net157 RN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X36 VDD net146 s VDD LPPFET W=0.66U L=0.12U M=1 
X37 s net146 VSS VSS LPNFET W=0.44U L=0.12U M=1 
X38 VDD net151 QN VDD LPPFET W=2.4U L=0.12U M=1 
X39 QN net151 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X4 pm c nminsi VDD LPPFET W=0.28U L=0.12U M=1 
X40 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X41 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X42 VDD CK cn VDD LPPFET W=0.44U L=0.12U M=1 
X43 cn CK VSS VSS LPNFET W=0.32U L=0.12U M=1 
X5 m SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X6 m pm net94 VDD LPPFET W=0.46U L=0.12U M=1 
X7 net94 net157 VDD VDD LPPFET W=0.62U L=0.12U M=1 
X8 net146 SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X9 net104 s net94 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS SDFFSRX4TS 

**** 
*.SUBCKT SDFFSRXLTS Q QN CK D RN SE SI SN 
.SUBCKT SDFFSRXLTS Q QN CK D RN SE SI SN VSS VDD
X0 VDD D hnet32 VDD LPPFET W=0.28U L=0.12U M=1 
X1 hnet32 SE nminsi VDD LPPFET W=0.28U L=0.12U M=1 
X10 net146 c net104 VDD LPPFET W=0.28U L=0.12U M=1 
X11 net146 cn m VDD LPPFET W=0.28U L=0.12U M=1 
X12 net115 D VSS VSS LPNFET W=0.2U L=0.12U M=1 
X13 nminsi nmse net115 VSS LPNFET W=0.2U L=0.12U M=1 
X14 net121 SI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X15 nminsi SE net121 VSS LPNFET W=0.2U L=0.12U M=1 
X16 pm cn nminsi VSS LPNFET W=0.2U L=0.12U M=1 
X17 m net157 net140 VSS LPNFET W=0.2U L=0.12U M=1 
X18 m pm net140 VSS LPNFET W=0.3U L=0.12U M=1 
X19 net146 net157 net140 VSS LPNFET W=0.2U L=0.12U M=1 
X2 VDD SI hnet36 VDD LPPFET W=0.28U L=0.12U M=1 
X20 net137 s net140 VSS LPNFET W=0.2U L=0.12U M=1 
X21 net140 SN VSS VSS LPNFET W=0.4U L=0.12U M=1 
X22 net146 cn net137 VSS LPNFET W=0.2U L=0.12U M=1 
X23 net146 c m VSS LPNFET W=0.2U L=0.12U M=1 
X24 hnet38 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X25 pm c hnet38 VSS LPNFET W=0.2U L=0.12U M=1 
X26 hnet40 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X27 VDD m hnet40 VDD LPPFET W=0.28U L=0.12U M=1 
X28 VDD s net151 VDD LPPFET W=0.28U L=0.12U M=1 
X29 net151 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 hnet36 nmse nminsi VDD LPPFET W=0.28U L=0.12U M=1 
X30 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X31 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X32 VDD s Q VDD LPPFET W=0.34U L=0.12U M=1 
X33 Q s VSS VSS LPNFET W=0.24U L=0.12U M=1 
X34 VDD RN net157 VDD LPPFET W=0.28U L=0.12U M=1 
X35 net157 RN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X36 VDD net146 s VDD LPPFET W=0.28U L=0.12U M=1 
X37 s net146 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X38 VDD net151 QN VDD LPPFET W=0.34U L=0.12U M=1 
X39 QN net151 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X4 pm c nminsi VDD LPPFET W=0.28U L=0.12U M=1 
X40 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X41 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X42 VDD CK cn VDD LPPFET W=0.42U L=0.12U M=1 
X43 cn CK VSS VSS LPNFET W=0.3U L=0.12U M=1 
X5 m SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X6 m pm net94 VDD LPPFET W=0.42U L=0.12U M=1 
X7 net94 net157 VDD VDD LPPFET W=0.56U L=0.12U M=1 
X8 net146 SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X9 net104 s net94 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS SDFFSRXLTS 

**** 
*.SUBCKT SDFFSX1TS Q QN CK D SE SI SN 
.SUBCKT SDFFSX1TS Q QN CK D SE SI SN VSS VDD
X0 VDD D hnet29 VDD LPPFET W=0.28U L=0.12U M=1 
X1 hnet29 SE nminsi VDD LPPFET W=0.28U L=0.12U M=1 
X10 net128 cn m VDD LPPFET W=0.28U L=0.12U M=1 
X11 net101 D VSS VSS LPNFET W=0.2U L=0.12U M=1 
X12 nminsi nmse net101 VSS LPNFET W=0.2U L=0.12U M=1 
X13 net109 SI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X14 nminsi SE net109 VSS LPNFET W=0.2U L=0.12U M=1 
X15 pm cn nminsi VSS LPNFET W=0.2U L=0.12U M=1 
X16 m pm net122 VSS LPNFET W=0.3U L=0.12U M=1 
X17 net119 s net122 VSS LPNFET W=0.2U L=0.12U M=1 
X18 net122 SN VSS VSS LPNFET W=0.4U L=0.12U M=1 
X19 net128 cn net119 VSS LPNFET W=0.2U L=0.12U M=1 
X2 VDD SI hnet33 VDD LPPFET W=0.28U L=0.12U M=1 
X20 net128 c m VSS LPNFET W=0.2U L=0.12U M=1 
X21 hnet35 m VSS VSS LPNFET W=0.22U L=0.12U M=1 
X22 pm c hnet35 VSS LPNFET W=0.22U L=0.12U M=1 
X23 hnet37 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X24 VDD m hnet37 VDD LPPFET W=0.28U L=0.12U M=1 
X25 VDD s net133 VDD LPPFET W=0.28U L=0.12U M=1 
X26 net133 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X27 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X28 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X29 VDD s Q VDD LPPFET W=0.64U L=0.12U M=1 
X3 hnet33 nmse nminsi VDD LPPFET W=0.28U L=0.12U M=1 
X30 Q s VSS VSS LPNFET W=0.46U L=0.12U M=1 
X31 VDD net128 s VDD LPPFET W=0.28U L=0.12U M=1 
X32 s net128 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X33 VDD net133 QN VDD LPPFET W=0.64U L=0.12U M=1 
X34 QN net133 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X35 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X36 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X37 VDD CK cn VDD LPPFET W=0.34U L=0.12U M=1 
X38 cn CK VSS VSS LPNFET W=0.24U L=0.12U M=1 
X4 pm c nminsi VDD LPPFET W=0.28U L=0.12U M=1 
X5 net83 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X6 m SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X7 m pm VDD VDD LPPFET W=0.28U L=0.12U M=1 
X8 net128 SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X9 net128 c net83 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS SDFFSX1TS 

**** 
*.SUBCKT SDFFSX2TS Q QN CK D SE SI SN 
.SUBCKT SDFFSX2TS Q QN CK D SE SI SN VSS VDD
X0 VDD D hnet29 VDD LPPFET W=0.28U L=0.12U M=1 
X1 hnet29 SE nminsi VDD LPPFET W=0.28U L=0.12U M=1 
X10 net128 cn m VDD LPPFET W=0.28U L=0.12U M=1 
X11 net103 D VSS VSS LPNFET W=0.2U L=0.12U M=1 
X12 nminsi nmse net103 VSS LPNFET W=0.2U L=0.12U M=1 
X13 net109 SI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X14 nminsi SE net109 VSS LPNFET W=0.2U L=0.12U M=1 
X15 pm cn nminsi VSS LPNFET W=0.22U L=0.12U M=1 
X16 m pm net122 VSS LPNFET W=0.3U L=0.12U M=1 
X17 net119 s net122 VSS LPNFET W=0.2U L=0.12U M=1 
X18 net122 SN VSS VSS LPNFET W=0.4U L=0.12U M=1 
X19 net128 cn net119 VSS LPNFET W=0.2U L=0.12U M=1 
X2 VDD SI hnet33 VDD LPPFET W=0.28U L=0.12U M=1 
X20 net128 c m VSS LPNFET W=0.2U L=0.12U M=1 
X21 hnet35 m VSS VSS LPNFET W=0.22U L=0.12U M=1 
X22 pm c hnet35 VSS LPNFET W=0.22U L=0.12U M=1 
X23 hnet37 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X24 VDD m hnet37 VDD LPPFET W=0.28U L=0.12U M=1 
X25 VDD s net133 VDD LPPFET W=0.3U L=0.12U M=1 
X26 net133 s VSS VSS LPNFET W=0.22U L=0.12U M=1 
X27 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X28 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X29 VDD s Q VDD LPPFET W=1.28U L=0.12U M=1 
X3 hnet33 nmse nminsi VDD LPPFET W=0.28U L=0.12U M=1 
X30 Q s VSS VSS LPNFET W=0.92U L=0.12U M=1 
X31 VDD net128 s VDD LPPFET W=0.36U L=0.12U M=1 
X32 s net128 VSS VSS LPNFET W=0.26U L=0.12U M=1 
X33 VDD net133 QN VDD LPPFET W=1.28U L=0.12U M=1 
X34 QN net133 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X35 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X36 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X37 VDD CK cn VDD LPPFET W=0.42U L=0.12U M=1 
X38 cn CK VSS VSS LPNFET W=0.3U L=0.12U M=1 
X4 pm c nminsi VDD LPPFET W=0.28U L=0.12U M=1 
X5 net94 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X6 m SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X7 m pm VDD VDD LPPFET W=0.28U L=0.12U M=1 
X8 net128 SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X9 net128 c net94 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS SDFFSX2TS 

**** 
*.SUBCKT SDFFSX4TS Q QN CK D SE SI SN 
.SUBCKT SDFFSX4TS Q QN CK D SE SI SN VSS VDD
X0 VDD D hnet29 VDD LPPFET W=0.28U L=0.12U M=1 
X1 hnet29 SE nminsi VDD LPPFET W=0.28U L=0.12U M=1 
X10 net128 cn m VDD LPPFET W=0.28U L=0.12U M=1 
X11 net103 D VSS VSS LPNFET W=0.2U L=0.12U M=1 
X12 nminsi nmse net103 VSS LPNFET W=0.2U L=0.12U M=1 
X13 net109 SI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X14 nminsi SE net109 VSS LPNFET W=0.2U L=0.12U M=1 
X15 pm cn nminsi VSS LPNFET W=0.2U L=0.12U M=1 
X16 m pm net122 VSS LPNFET W=0.34U L=0.12U M=1 
X17 net119 s net122 VSS LPNFET W=0.2U L=0.12U M=1 
X18 net122 SN VSS VSS LPNFET W=0.46U L=0.12U M=1 
X19 net128 cn net119 VSS LPNFET W=0.2U L=0.12U M=1 
X2 VDD SI hnet33 VDD LPPFET W=0.28U L=0.12U M=1 
X20 net128 c m VSS LPNFET W=0.22U L=0.12U M=1 
X21 hnet35 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X22 pm c hnet35 VSS LPNFET W=0.2U L=0.12U M=1 
X23 hnet37 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X24 VDD m hnet37 VDD LPPFET W=0.28U L=0.12U M=1 
X25 VDD s net133 VDD LPPFET W=0.62U L=0.12U M=1 
X26 net133 s VSS VSS LPNFET W=0.44U L=0.12U M=1 
X27 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X28 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X29 VDD s Q VDD LPPFET W=2.56U L=0.12U M=1 
X3 hnet33 nmse nminsi VDD LPPFET W=0.28U L=0.12U M=1 
X30 Q s VSS VSS LPNFET W=1.84U L=0.12U M=1 
X31 VDD net128 s VDD LPPFET W=0.66U L=0.12U M=1 
X32 s net128 VSS VSS LPNFET W=0.48U L=0.12U M=1 
X33 VDD net133 QN VDD LPPFET W=2.56U L=0.12U M=1 
X34 QN net133 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X35 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X36 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X37 VDD CK cn VDD LPPFET W=0.42U L=0.12U M=1 
X38 cn CK VSS VSS LPNFET W=0.3U L=0.12U M=1 
X4 pm c nminsi VDD LPPFET W=0.28U L=0.12U M=1 
X5 net94 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X6 m SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X7 m pm VDD VDD LPPFET W=0.28U L=0.12U M=1 
X8 net128 SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X9 net128 c net94 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS SDFFSX4TS 

**** 
*.SUBCKT SDFFSXLTS Q QN CK D SE SI SN 
.SUBCKT SDFFSXLTS Q QN CK D SE SI SN VSS VDD
X0 VDD D hnet29 VDD LPPFET W=0.28U L=0.12U M=1 
X1 hnet29 SE nminsi VDD LPPFET W=0.28U L=0.12U M=1 
X10 net128 cn m VDD LPPFET W=0.28U L=0.12U M=1 
X11 net101 D VSS VSS LPNFET W=0.2U L=0.12U M=1 
X12 nminsi nmse net101 VSS LPNFET W=0.2U L=0.12U M=1 
X13 net109 SI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X14 nminsi SE net109 VSS LPNFET W=0.2U L=0.12U M=1 
X15 pm cn nminsi VSS LPNFET W=0.2U L=0.12U M=1 
X16 m pm net122 VSS LPNFET W=0.3U L=0.12U M=1 
X17 net119 s net122 VSS LPNFET W=0.2U L=0.12U M=1 
X18 net122 SN VSS VSS LPNFET W=0.4U L=0.12U M=1 
X19 net128 cn net119 VSS LPNFET W=0.2U L=0.12U M=1 
X2 VDD SI hnet33 VDD LPPFET W=0.28U L=0.12U M=1 
X20 net128 c m VSS LPNFET W=0.2U L=0.12U M=1 
X21 hnet35 m VSS VSS LPNFET W=0.22U L=0.12U M=1 
X22 pm c hnet35 VSS LPNFET W=0.22U L=0.12U M=1 
X23 hnet37 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X24 VDD m hnet37 VDD LPPFET W=0.28U L=0.12U M=1 
X25 VDD s net133 VDD LPPFET W=0.28U L=0.12U M=1 
X26 net133 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X27 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X28 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X29 VDD s Q VDD LPPFET W=0.34U L=0.12U M=1 
X3 hnet33 nmse nminsi VDD LPPFET W=0.28U L=0.12U M=1 
X30 Q s VSS VSS LPNFET W=0.24U L=0.12U M=1 
X31 VDD net128 s VDD LPPFET W=0.28U L=0.12U M=1 
X32 s net128 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X33 VDD net133 QN VDD LPPFET W=0.34U L=0.12U M=1 
X34 QN net133 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X35 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X36 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X37 VDD CK cn VDD LPPFET W=0.34U L=0.12U M=1 
X38 cn CK VSS VSS LPNFET W=0.24U L=0.12U M=1 
X4 pm c nminsi VDD LPPFET W=0.28U L=0.12U M=1 
X5 net83 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X6 m SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X7 m pm VDD VDD LPPFET W=0.28U L=0.12U M=1 
X8 net128 SN VDD VDD LPPFET W=0.28U L=0.12U M=1 
X9 net128 c net83 VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS SDFFSXLTS 

**** 
*.SUBCKT SDFFTRX1TS Q QN CK D RN SE SI 
.SUBCKT SDFFTRX1TS Q QN CK D RN SE SI VSS VDD
X0 VDD SE hnet29 VDD LPPFET W=0.28U L=0.12U M=1 
X1 hnet29 RN net99 VDD LPPFET W=0.28U L=0.12U M=1 
X10 pm c net99 VDD LPPFET W=0.28U L=0.12U M=1 
X11 net117 c net87 VDD LPPFET W=0.28U L=0.12U M=1 
X12 net87 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X13 net117 cn m VDD LPPFET W=0.28U L=0.12U M=1 
X14 net93 RN VSS VSS LPNFET W=0.28U L=0.12U M=1 
X15 net98 D net93 VSS LPNFET W=0.28U L=0.12U M=1 
X16 net99 nmse net98 VSS LPNFET W=0.28U L=0.12U M=1 
X17 net104 SI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X18 net99 SE net104 VSS LPNFET W=0.2U L=0.12U M=1 
X19 pm cn net99 VSS LPNFET W=0.2U L=0.12U M=1 
X2 VDD D hnet33 VDD LPPFET W=0.36U L=0.12U M=1 
X20 net117 cn net114 VSS LPNFET W=0.2U L=0.12U M=1 
X21 net114 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X22 net117 c m VSS LPNFET W=0.2U L=0.12U M=1 
X23 VDD s net118 VDD LPPFET W=0.28U L=0.12U M=1 
X24 net118 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X25 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X26 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X27 VDD net117 s VDD LPPFET W=0.28U L=0.12U M=1 
X28 s net117 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X29 VDD pm m VDD LPPFET W=0.28U L=0.12U M=1 
X3 hnet33 SE net99 VDD LPPFET W=0.36U L=0.12U M=1 
X30 m pm VSS VSS LPNFET W=0.2U L=0.12U M=1 
X31 VDD s Q VDD LPPFET W=0.64U L=0.12U M=1 
X32 Q s VSS VSS LPNFET W=0.46U L=0.12U M=1 
X33 VDD net118 QN VDD LPPFET W=0.64U L=0.12U M=1 
X34 QN net118 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X35 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X36 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X37 VDD CK cn VDD LPPFET W=0.42U L=0.12U M=1 
X38 cn CK VSS VSS LPNFET W=0.3U L=0.12U M=1 
X4 VDD SI hnet37 VDD LPPFET W=0.28U L=0.12U M=1 
X5 hnet37 nmse net99 VDD LPPFET W=0.28U L=0.12U M=1 
X6 VDD m hnet41 VDD LPPFET W=0.28U L=0.12U M=1 
X7 hnet41 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X8 hnet45 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X9 pm c hnet45 VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS SDFFTRX1TS 

**** 
*.SUBCKT SDFFTRX2TS Q QN CK D RN SE SI 
.SUBCKT SDFFTRX2TS Q QN CK D RN SE SI VSS VDD
X0 VDD SE hnet29 VDD LPPFET W=0.28U L=0.12U M=1 
X1 hnet29 RN net99 VDD LPPFET W=0.28U L=0.12U M=1 
X10 pm c net99 VDD LPPFET W=0.28U L=0.12U M=1 
X11 net117 c net87 VDD LPPFET W=0.28U L=0.12U M=1 
X12 net87 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X13 net117 cn m VDD LPPFET W=0.28U L=0.12U M=1 
X14 net93 RN VSS VSS LPNFET W=0.28U L=0.12U M=1 
X15 net98 D net93 VSS LPNFET W=0.28U L=0.12U M=1 
X16 net99 nmse net98 VSS LPNFET W=0.28U L=0.12U M=1 
X17 net104 SI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X18 net99 SE net104 VSS LPNFET W=0.2U L=0.12U M=1 
X19 pm cn net99 VSS LPNFET W=0.2U L=0.12U M=1 
X2 VDD D hnet33 VDD LPPFET W=0.36U L=0.12U M=1 
X20 net117 cn net114 VSS LPNFET W=0.2U L=0.12U M=1 
X21 net114 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X22 net117 c m VSS LPNFET W=0.2U L=0.12U M=1 
X23 VDD s net118 VDD LPPFET W=0.3U L=0.12U M=1 
X24 net118 s VSS VSS LPNFET W=0.22U L=0.12U M=1 
X25 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X26 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X27 VDD net117 s VDD LPPFET W=0.36U L=0.12U M=1 
X28 s net117 VSS VSS LPNFET W=0.26U L=0.12U M=1 
X29 VDD pm m VDD LPPFET W=0.28U L=0.12U M=1 
X3 hnet33 SE net99 VDD LPPFET W=0.36U L=0.12U M=1 
X30 m pm VSS VSS LPNFET W=0.2U L=0.12U M=1 
X31 VDD s Q VDD LPPFET W=1.28U L=0.12U M=1 
X32 Q s VSS VSS LPNFET W=0.92U L=0.12U M=1 
X33 VDD net118 QN VDD LPPFET W=1.28U L=0.12U M=1 
X34 QN net118 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X35 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X36 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X37 VDD CK cn VDD LPPFET W=0.42U L=0.12U M=1 
X38 cn CK VSS VSS LPNFET W=0.3U L=0.12U M=1 
X4 VDD SI hnet37 VDD LPPFET W=0.28U L=0.12U M=1 
X5 hnet37 nmse net99 VDD LPPFET W=0.28U L=0.12U M=1 
X6 VDD m hnet41 VDD LPPFET W=0.28U L=0.12U M=1 
X7 hnet41 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X8 hnet45 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X9 pm c hnet45 VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS SDFFTRX2TS 

**** 
*.SUBCKT SDFFTRX4TS Q QN CK D RN SE SI 
.SUBCKT SDFFTRX4TS Q QN CK D RN SE SI VSS VDD
X0 VDD SE hnet29 VDD LPPFET W=0.28U L=0.12U M=1 
X1 hnet29 RN net99 VDD LPPFET W=0.28U L=0.12U M=1 
X10 pm c net99 VDD LPPFET W=0.28U L=0.12U M=1 
X11 net117 c net87 VDD LPPFET W=0.28U L=0.12U M=1 
X12 net87 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X13 net117 cn m VDD LPPFET W=0.28U L=0.12U M=1 
X14 net93 RN VSS VSS LPNFET W=0.28U L=0.12U M=1 
X15 net98 D net93 VSS LPNFET W=0.28U L=0.12U M=1 
X16 net99 nmse net98 VSS LPNFET W=0.28U L=0.12U M=1 
X17 net104 SI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X18 net99 SE net104 VSS LPNFET W=0.2U L=0.12U M=1 
X19 pm cn net99 VSS LPNFET W=0.2U L=0.12U M=1 
X2 VDD D hnet33 VDD LPPFET W=0.36U L=0.12U M=1 
X20 net117 cn net114 VSS LPNFET W=0.2U L=0.12U M=1 
X21 net114 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X22 net117 c m VSS LPNFET W=0.22U L=0.12U M=1 
X23 VDD s net118 VDD LPPFET W=0.62U L=0.12U M=1 
X24 net118 s VSS VSS LPNFET W=0.4U L=0.12U M=1 
X25 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X26 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X27 VDD net117 s VDD LPPFET W=0.66U L=0.12U M=1 
X28 s net117 VSS VSS LPNFET W=0.44U L=0.12U M=1 
X29 VDD pm m VDD LPPFET W=0.28U L=0.12U M=1 
X3 hnet33 SE net99 VDD LPPFET W=0.36U L=0.12U M=1 
X30 m pm VSS VSS LPNFET W=0.22U L=0.12U M=1 
X31 VDD s Q VDD LPPFET W=2.4U L=0.12U M=1 
X32 Q s VSS VSS LPNFET W=1.84U L=0.12U M=1 
X33 VDD net118 QN VDD LPPFET W=2.4U L=0.12U M=1 
X34 QN net118 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X35 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X36 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X37 VDD CK cn VDD LPPFET W=0.44U L=0.12U M=1 
X38 cn CK VSS VSS LPNFET W=0.32U L=0.12U M=1 
X4 VDD SI hnet37 VDD LPPFET W=0.28U L=0.12U M=1 
X5 hnet37 nmse net99 VDD LPPFET W=0.28U L=0.12U M=1 
X6 VDD m hnet41 VDD LPPFET W=0.28U L=0.12U M=1 
X7 hnet41 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X8 hnet45 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X9 pm c hnet45 VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS SDFFTRX4TS 

**** 
*.SUBCKT SDFFTRXLTS Q QN CK D RN SE SI 
.SUBCKT SDFFTRXLTS Q QN CK D RN SE SI VSS VDD
X0 VDD SE hnet29 VDD LPPFET W=0.28U L=0.12U M=1 
X1 hnet29 RN net99 VDD LPPFET W=0.28U L=0.12U M=1 
X10 pm c net99 VDD LPPFET W=0.28U L=0.12U M=1 
X11 net117 c net87 VDD LPPFET W=0.28U L=0.12U M=1 
X12 net87 s VDD VDD LPPFET W=0.28U L=0.12U M=1 
X13 net117 cn m VDD LPPFET W=0.28U L=0.12U M=1 
X14 net93 RN VSS VSS LPNFET W=0.28U L=0.12U M=1 
X15 net98 D net93 VSS LPNFET W=0.28U L=0.12U M=1 
X16 net99 nmse net98 VSS LPNFET W=0.28U L=0.12U M=1 
X17 net104 SI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X18 net99 SE net104 VSS LPNFET W=0.2U L=0.12U M=1 
X19 pm cn net99 VSS LPNFET W=0.2U L=0.12U M=1 
X2 VDD D hnet33 VDD LPPFET W=0.36U L=0.12U M=1 
X20 net117 cn net114 VSS LPNFET W=0.2U L=0.12U M=1 
X21 net114 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X22 net117 c m VSS LPNFET W=0.2U L=0.12U M=1 
X23 VDD s net118 VDD LPPFET W=0.28U L=0.12U M=1 
X24 net118 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X25 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X26 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X27 VDD net117 s VDD LPPFET W=0.28U L=0.12U M=1 
X28 s net117 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X29 VDD pm m VDD LPPFET W=0.28U L=0.12U M=1 
X3 hnet33 SE net99 VDD LPPFET W=0.36U L=0.12U M=1 
X30 m pm VSS VSS LPNFET W=0.2U L=0.12U M=1 
X31 VDD s Q VDD LPPFET W=0.34U L=0.12U M=1 
X32 Q s VSS VSS LPNFET W=0.24U L=0.12U M=1 
X33 VDD net118 QN VDD LPPFET W=0.34U L=0.12U M=1 
X34 QN net118 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X35 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X36 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X37 VDD CK cn VDD LPPFET W=0.42U L=0.12U M=1 
X38 cn CK VSS VSS LPNFET W=0.3U L=0.12U M=1 
X4 VDD SI hnet37 VDD LPPFET W=0.28U L=0.12U M=1 
X5 hnet37 nmse net99 VDD LPPFET W=0.28U L=0.12U M=1 
X6 VDD m hnet41 VDD LPPFET W=0.28U L=0.12U M=1 
X7 hnet41 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X8 hnet45 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X9 pm c hnet45 VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS SDFFTRXLTS 

**** 
*.SUBCKT SDFFX1TS Q QN CK D SE SI 
.SUBCKT SDFFX1TS Q QN CK D SE SI VSS VDD
X0 VDD SE hnet26 VDD LPPFET W=0.28U L=0.12U M=1 
X1 hnet26 D net50 VDD LPPFET W=0.28U L=0.12U M=1 
X10 hnet28 m VSS VSS LPNFET W=0.58U L=0.12U M=1 
X11 net82 c hnet28 VSS LPNFET W=0.58U L=0.12U M=1 
X12 hnet30 cn net82 VDD LPPFET W=0.8U L=0.12U M=1 
X13 VDD m hnet30 VDD LPPFET W=0.8U L=0.12U M=1 
X14 hnet34 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X15 net82 cn hnet34 VSS LPNFET W=0.2U L=0.12U M=1 
X16 hnet36 c net82 VDD LPPFET W=0.28U L=0.12U M=1 
X17 VDD s hnet36 VDD LPPFET W=0.28U L=0.12U M=1 
X18 hnet40 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X19 pm c hnet40 VSS LPNFET W=0.2U L=0.12U M=1 
X2 net58 SE net67 VSS LPNFET W=0.2U L=0.12U M=1 
X20 hnet42 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X21 VDD m hnet42 VDD LPPFET W=0.28U L=0.12U M=1 
X22 VDD s QN VDD LPPFET W=0.64U L=0.12U M=1 
X23 QN s VSS VSS LPNFET W=0.46U L=0.12U M=1 
X24 VDD net82 s VDD LPPFET W=0.36U L=0.12U M=1 
X25 s net82 VSS VSS LPNFET W=0.26U L=0.12U M=1 
X26 VDD pm m VDD LPPFET W=0.3U L=0.12U M=1 
X27 m pm VSS VSS LPNFET W=0.2U L=0.12U M=1 
X28 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X29 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 net58 D net61 VSS LPNFET W=0.2U L=0.12U M=1 
X30 VDD cn c VDD LPPFET W=0.3U L=0.12U M=1 
X31 c cn VSS VSS LPNFET W=0.22U L=0.12U M=1 
X32 VDD CK cn VDD LPPFET W=0.46U L=0.12U M=1 
X33 cn CK VSS VSS LPNFET W=0.34U L=0.12U M=1 
X34 VDD net82 Q VDD LPPFET W=0.64U L=0.12U M=1 
X35 Q net82 VSS VSS LPNFET W=0.42U L=0.12U M=1 
X4 net61 nmse VSS VSS LPNFET W=0.2U L=0.12U M=1 
X5 pm cn net58 VSS LPNFET W=0.2U L=0.12U M=1 
X6 net67 SI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X7 net50 nmse net76 VDD LPPFET W=0.28U L=0.12U M=1 
X8 pm c net50 VDD LPPFET W=0.28U L=0.12U M=1 
X9 net76 SI VDD VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS SDFFX1TS 

**** 
*.SUBCKT SDFFX2TS Q QN CK D SE SI 
.SUBCKT SDFFX2TS Q QN CK D SE SI VSS VDD
X0 VDD SE hnet26 VDD LPPFET W=0.32U L=0.12U M=1 
X1 hnet26 D net50 VDD LPPFET W=0.32U L=0.12U M=1 
X10 hnet28 m VSS VSS LPNFET W=0.92U L=0.12U M=1 
X11 net82 c hnet28 VSS LPNFET W=0.92U L=0.12U M=1 
X12 hnet30 cn net82 VDD LPPFET W=1.3U L=0.12U M=1 
X13 VDD m hnet30 VDD LPPFET W=1.3U L=0.12U M=1 
X14 hnet34 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X15 net82 cn hnet34 VSS LPNFET W=0.2U L=0.12U M=1 
X16 hnet36 c net82 VDD LPPFET W=0.26U L=0.12U M=1 
X17 VDD s hnet36 VDD LPPFET W=0.26U L=0.12U M=1 
X18 hnet40 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X19 pm c hnet40 VSS LPNFET W=0.2U L=0.12U M=1 
X2 net58 SE net67 VSS LPNFET W=0.2U L=0.12U M=1 
X20 hnet42 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X21 VDD m hnet42 VDD LPPFET W=0.28U L=0.12U M=1 
X22 VDD s QN VDD LPPFET W=1.3U L=0.12U M=1 
X23 QN s VSS VSS LPNFET W=0.92U L=0.12U M=1 
X24 VDD net82 s VDD LPPFET W=0.62U L=0.12U M=1 
X25 s net82 VSS VSS LPNFET W=0.44U L=0.12U M=1 
X26 VDD pm m VDD LPPFET W=0.44U L=0.12U M=1 
X27 m pm VSS VSS LPNFET W=0.36U L=0.12U M=1 
X28 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X29 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 net58 D net61 VSS LPNFET W=0.22U L=0.12U M=1 
X30 VDD cn c VDD LPPFET W=0.44U L=0.12U M=1 
X31 c cn VSS VSS LPNFET W=0.3U L=0.12U M=1 
X32 VDD CK cn VDD LPPFET W=0.66U L=0.12U M=1 
X33 cn CK VSS VSS LPNFET W=0.48U L=0.12U M=1 
X34 VDD net82 Q VDD LPPFET W=1.28U L=0.12U M=1 
X35 Q net82 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X4 net61 nmse VSS VSS LPNFET W=0.22U L=0.12U M=1 
X5 pm cn net58 VSS LPNFET W=0.22U L=0.12U M=1 
X6 net67 SI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X7 net50 nmse net76 VDD LPPFET W=0.28U L=0.12U M=1 
X8 pm c net50 VDD LPPFET W=0.32U L=0.12U M=1 
X9 net76 SI VDD VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS SDFFX2TS 

**** 
*.SUBCKT SDFFX4TS Q QN CK D SE SI 
.SUBCKT SDFFX4TS Q QN CK D SE SI VSS VDD
X0 VDD SE hnet26 VDD LPPFET W=0.58U L=0.12U M=1 
X1 hnet26 D net50 VDD LPPFET W=0.58U L=0.12U M=1 
X10 hnet28 cn net82 VDD LPPFET W=0.98U L=0.12U M=1 
X11 VDD m hnet30 VDD LPPFET W=0.98U L=0.12U M=1 
X12 VDD m hnet32 VDD LPPFET W=0.98U L=0.12U M=1 
X13 VDD m hnet28 VDD LPPFET W=0.98U L=0.12U M=1 
X14 net62 SE net71 VSS LPNFET W=0.2U L=0.12U M=1 
X15 net62 D net65 VSS LPNFET W=0.42U L=0.12U M=1 
X16 net65 nmse VSS VSS LPNFET W=0.42U L=0.12U M=1 
X17 pm cn net62 VSS LPNFET W=0.42U L=0.12U M=1 
X18 net71 SI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X19 net50 nmse net80 VDD LPPFET W=0.28U L=0.12U M=1 
X2 hnet29 m VSS VSS LPNFET W=0.66U L=0.12U M=1 
X20 pm c net50 VDD LPPFET W=0.58U L=0.12U M=1 
X21 net80 SI VDD VDD LPPFET W=0.28U L=0.12U M=1 
X22 hnet38 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X23 net82 cn hnet38 VSS LPNFET W=0.2U L=0.12U M=1 
X24 hnet40 c net82 VDD LPPFET W=0.28U L=0.12U M=1 
X25 VDD s hnet40 VDD LPPFET W=0.28U L=0.12U M=1 
X26 hnet44 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X27 pm c hnet44 VSS LPNFET W=0.2U L=0.12U M=1 
X28 hnet46 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X29 VDD m hnet46 VDD LPPFET W=0.28U L=0.12U M=1 
X3 hnet31 m VSS VSS LPNFET W=0.66U L=0.12U M=1 
X30 VDD s QN VDD LPPFET W=2.4U L=0.12U M=1 
X31 QN s VSS VSS LPNFET W=1.84U L=0.12U M=1 
X32 VDD net82 s VDD LPPFET W=1.14U L=0.12U M=1 
X33 s net82 VSS VSS LPNFET W=0.82U L=0.12U M=1 
X34 VDD pm m VDD LPPFET W=0.88U L=0.12U M=1 
X35 m pm VSS VSS LPNFET W=0.62U L=0.12U M=1 
X36 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X37 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X38 VDD cn c VDD LPPFET W=0.8U L=0.12U M=1 
X39 c cn VSS VSS LPNFET W=0.54U L=0.12U M=1 
X4 hnet35 m VSS VSS LPNFET W=0.66U L=0.12U M=1 
X40 VDD CK cn VDD LPPFET W=1.06U L=0.12U M=1 
X41 cn CK VSS VSS LPNFET W=0.7U L=0.12U M=1 
X42 VDD net82 Q VDD LPPFET W=2.4U L=0.12U M=1 
X43 Q net82 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X5 net82 c hnet29 VSS LPNFET W=0.66U L=0.12U M=1 
X6 net82 c hnet31 VSS LPNFET W=0.66U L=0.12U M=1 
X7 net82 c hnet35 VSS LPNFET W=0.66U L=0.12U M=1 
X8 hnet30 cn net82 VDD LPPFET W=0.98U L=0.12U M=1 
X9 hnet32 cn net82 VDD LPPFET W=0.98U L=0.12U M=1 
.ENDS SDFFX4TS 

**** 
*.SUBCKT SDFFXLTS Q QN CK D SE SI 
.SUBCKT SDFFXLTS Q QN CK D SE SI VSS VDD
X0 VDD SE hnet26 VDD LPPFET W=0.28U L=0.12U M=1 
X1 hnet26 D net50 VDD LPPFET W=0.28U L=0.12U M=1 
X10 hnet28 m VSS VSS LPNFET W=0.36U L=0.12U M=1 
X11 net82 c hnet28 VSS LPNFET W=0.36U L=0.12U M=1 
X12 hnet30 cn net82 VDD LPPFET W=0.5U L=0.12U M=1 
X13 VDD m hnet30 VDD LPPFET W=0.5U L=0.12U M=1 
X14 hnet34 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X15 net82 cn hnet34 VSS LPNFET W=0.2U L=0.12U M=1 
X16 hnet36 c net82 VDD LPPFET W=0.28U L=0.12U M=1 
X17 VDD s hnet36 VDD LPPFET W=0.28U L=0.12U M=1 
X18 hnet40 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X19 pm c hnet40 VSS LPNFET W=0.2U L=0.12U M=1 
X2 net58 SE net67 VSS LPNFET W=0.2U L=0.12U M=1 
X20 hnet42 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X21 VDD m hnet42 VDD LPPFET W=0.28U L=0.12U M=1 
X22 VDD s QN VDD LPPFET W=0.34U L=0.12U M=1 
X23 QN s VSS VSS LPNFET W=0.24U L=0.12U M=1 
X24 VDD net82 s VDD LPPFET W=0.28U L=0.12U M=1 
X25 s net82 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X26 VDD pm m VDD LPPFET W=0.28U L=0.12U M=1 
X27 m pm VSS VSS LPNFET W=0.2U L=0.12U M=1 
X28 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X29 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 net58 D net61 VSS LPNFET W=0.2U L=0.12U M=1 
X30 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X31 c cn VSS VSS LPNFET W=0.18U L=0.12U M=1 
X32 VDD CK cn VDD LPPFET W=0.38U L=0.12U M=1 
X33 cn CK VSS VSS LPNFET W=0.26U L=0.12U M=1 
X34 VDD net82 Q VDD LPPFET W=0.34U L=0.12U M=1 
X35 Q net82 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X4 net61 nmse VSS VSS LPNFET W=0.2U L=0.12U M=1 
X5 pm cn net58 VSS LPNFET W=0.2U L=0.12U M=1 
X6 net67 SI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X7 net50 nmse net76 VDD LPPFET W=0.28U L=0.12U M=1 
X8 pm c net50 VDD LPPFET W=0.28U L=0.12U M=1 
X9 net76 SI VDD VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS SDFFXLTS 

**** 
*.SUBCKT SEDFFHQX1TS Q CK D E SE SI 
.SUBCKT SEDFFHQX1TS Q CK D E SE SI VSS VDD
X0 nmen SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X1 nmen E VSS VSS LPNFET W=0.2U L=0.12U M=1 
X10 hnet41 cn VSS VSS LPNFET W=0.36U L=0.12U M=1 
X11 pm nmsi hnet41 VSS LPNFET W=0.36U L=0.12U M=1 
X12 net89 CK VDD VDD LPPFET W=0.7U L=0.12U M=1 
X13 cn c net89 VDD LPPFET W=0.52U L=0.12U M=1 
X14 nmsi net79 nmin VDD LPPFET W=0.34U L=0.12U M=1 
X15 net121 cn m VDD LPPFET W=0.82U L=0.12U M=1 
X16 cn CK VSS VSS LPNFET W=0.2U L=0.12U M=1 
X17 nmsi net128 nmin VSS LPNFET W=0.24U L=0.12U M=1 
X18 net121 c m VSS LPNFET W=0.42U L=0.12U M=1 
X19 hnet43 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 VDD SE hnet27 VDD LPPFET W=0.36U L=0.12U M=1 
X20 nmsi nmen hnet43 VSS LPNFET W=0.2U L=0.12U M=1 
X21 hnet45 net130 nmsi VDD LPPFET W=0.28U L=0.12U M=1 
X22 VDD s hnet45 VDD LPPFET W=0.28U L=0.12U M=1 
X23 hnet49 SI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X24 nmsi SE hnet49 VSS LPNFET W=0.2U L=0.12U M=1 
X25 hnet51 nmse nmsi VDD LPPFET W=0.28U L=0.12U M=1 
X26 VDD SI hnet51 VDD LPPFET W=0.28U L=0.12U M=1 
X27 hnet55 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X28 pm c hnet55 VSS LPNFET W=0.2U L=0.12U M=1 
X29 hnet57 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X3 hnet27 E nmen VDD LPPFET W=0.36U L=0.12U M=1 
X30 VDD m hnet57 VDD LPPFET W=0.28U L=0.12U M=1 
X31 hnet61 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X32 net121 cn hnet61 VSS LPNFET W=0.2U L=0.12U M=1 
X33 hnet63 c net121 VDD LPPFET W=0.28U L=0.12U M=1 
X34 VDD s hnet63 VDD LPPFET W=0.28U L=0.12U M=1 
X35 VDD D nmin VDD LPPFET W=0.34U L=0.12U M=1 
X36 nmin D VSS VSS LPNFET W=0.24U L=0.12U M=1 
X37 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X38 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X39 VDD net79 net128 VDD LPPFET W=0.28U L=0.12U M=1 
X4 hnet33 nmse VSS VSS LPNFET W=0.2U L=0.12U M=1 
X40 net128 net79 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X41 VDD nmen net130 VDD LPPFET W=0.28U L=0.12U M=1 
X42 net130 nmen VSS VSS LPNFET W=0.2U L=0.12U M=1 
X43 VDD pm m VDD LPPFET W=0.84U L=0.12U M=1 
X44 m pm VSS VSS LPNFET W=0.44U L=0.12U M=1 
X45 VDD net121 s VDD LPPFET W=0.28U L=0.12U M=1 
X46 s net121 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X47 VDD net121 Q VDD LPPFET W=0.74U L=0.12U M=1 
X48 Q net121 VSS VSS LPNFET W=0.44U L=0.12U M=1 
X49 VDD net140 c VDD LPPFET W=0.78U L=0.12U M=1 
X5 net79 E hnet33 VSS LPNFET W=0.2U L=0.12U M=1 
X50 c net140 VSS VSS LPNFET W=0.28U L=0.12U M=1 
X51 VDD CK net140 VDD LPPFET W=0.28U L=0.12U M=1 
X52 net140 CK VSS VSS LPNFET W=0.28U L=0.12U M=1 
X6 VDD nmse net79 VDD LPPFET W=0.28U L=0.12U M=1 
X7 VDD E net79 VDD LPPFET W=0.28U L=0.12U M=1 
X8 VDD c hnet37 VDD LPPFET W=0.5U L=0.12U M=1 
X9 hnet37 nmsi pm VDD LPPFET W=0.5U L=0.12U M=1 
.ENDS SEDFFHQX1TS 

**** 
*.SUBCKT SEDFFHQX2TS Q CK D E SE SI 
.SUBCKT SEDFFHQX2TS Q CK D E SE SI VSS VDD
X0 nmen SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X1 nmen E VSS VSS LPNFET W=0.2U L=0.12U M=1 
X10 hnet41 cn VSS VSS LPNFET W=0.68U L=0.12U M=1 
X11 pm nmsi hnet41 VSS LPNFET W=0.68U L=0.12U M=1 
X12 net89 CK VDD VDD LPPFET W=0.9U L=0.12U M=1 
X13 cn c net89 VDD LPPFET W=0.68U L=0.12U M=1 
X14 nmsi net79 nmin VDD LPPFET W=0.64U L=0.12U M=1 
X15 net121 cn m VDD LPPFET W=1.38U L=0.12U M=1 
X16 cn CK VSS VSS LPNFET W=0.28U L=0.12U M=1 
X17 nmsi net128 nmin VSS LPNFET W=0.46U L=0.12U M=1 
X18 net121 c m VSS LPNFET W=0.68U L=0.12U M=1 
X19 hnet43 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 VDD SE hnet27 VDD LPPFET W=0.36U L=0.12U M=1 
X20 nmsi nmen hnet43 VSS LPNFET W=0.2U L=0.12U M=1 
X21 hnet45 net130 nmsi VDD LPPFET W=0.28U L=0.12U M=1 
X22 VDD s hnet45 VDD LPPFET W=0.28U L=0.12U M=1 
X23 hnet49 SI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X24 nmsi SE hnet49 VSS LPNFET W=0.2U L=0.12U M=1 
X25 hnet51 nmse nmsi VDD LPPFET W=0.28U L=0.12U M=1 
X26 VDD SI hnet51 VDD LPPFET W=0.28U L=0.12U M=1 
X27 hnet55 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X28 pm c hnet55 VSS LPNFET W=0.2U L=0.12U M=1 
X29 hnet57 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X3 hnet27 E nmen VDD LPPFET W=0.36U L=0.12U M=1 
X30 VDD m hnet57 VDD LPPFET W=0.28U L=0.12U M=1 
X31 hnet61 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X32 net121 cn hnet61 VSS LPNFET W=0.2U L=0.12U M=1 
X33 hnet63 c net121 VDD LPPFET W=0.28U L=0.12U M=1 
X34 VDD s hnet63 VDD LPPFET W=0.28U L=0.12U M=1 
X35 VDD D nmin VDD LPPFET W=0.64U L=0.12U M=1 
X36 nmin D VSS VSS LPNFET W=0.46U L=0.12U M=1 
X37 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X38 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X39 VDD net79 net128 VDD LPPFET W=0.28U L=0.12U M=1 
X4 hnet33 nmse VSS VSS LPNFET W=0.2U L=0.12U M=1 
X40 net128 net79 VSS VSS LPNFET W=0.18U L=0.12U M=1 
X41 VDD nmen net130 VDD LPPFET W=0.28U L=0.12U M=1 
X42 net130 nmen VSS VSS LPNFET W=0.2U L=0.12U M=1 
X43 VDD pm m VDD LPPFET W=1.38U L=0.12U M=1 
X44 m pm VSS VSS LPNFET W=0.68U L=0.12U M=1 
X45 VDD net121 s VDD LPPFET W=0.28U L=0.12U M=1 
X46 s net121 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X47 VDD net121 Q VDD LPPFET W=1.48U L=0.12U M=1 
X48 Q net121 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X49 VDD net140 c VDD LPPFET W=1.18U L=0.12U M=1 
X5 net79 E hnet33 VSS LPNFET W=0.2U L=0.12U M=1 
X50 c net140 VSS VSS LPNFET W=0.42U L=0.12U M=1 
X51 VDD CK net140 VDD LPPFET W=0.32U L=0.12U M=1 
X52 net140 CK VSS VSS LPNFET W=0.32U L=0.12U M=1 
X6 VDD nmse net79 VDD LPPFET W=0.28U L=0.12U M=1 
X7 VDD E net79 VDD LPPFET W=0.28U L=0.12U M=1 
X8 VDD c hnet37 VDD LPPFET W=0.94U L=0.12U M=1 
X9 hnet37 nmsi pm VDD LPPFET W=0.94U L=0.12U M=1 
.ENDS SEDFFHQX2TS 

**** 
*.SUBCKT SEDFFHQX4TS Q CK D E SE SI 
.SUBCKT SEDFFHQX4TS Q CK D E SE SI VSS VDD
X0 VDD c hnet31 VDD LPPFET W=0.86U L=0.12U M=1 
X1 hnet31 nmsi pm VDD LPPFET W=0.86U L=0.12U M=1 
X10 VDD SE hnet38 VDD LPPFET W=0.4U L=0.12U M=1 
X11 hnet38 E nmen VDD LPPFET W=0.4U L=0.12U M=1 
X12 hnet44 nmse VSS VSS LPNFET W=0.2U L=0.12U M=1 
X13 net86 E hnet44 VSS LPNFET W=0.2U L=0.12U M=1 
X14 VDD nmse net86 VDD LPPFET W=0.28U L=0.12U M=1 
X15 VDD E net86 VDD LPPFET W=0.28U L=0.12U M=1 
X16 cn c net89 VDD LPPFET W=0.62U L=0.12U M=1 
X17 net89 CK VDD VDD LPPFET W=0.84U L=0.12U M=1 
X18 net98 CK VDD VDD LPPFET W=0.72U L=0.12U M=1 
X19 cn c net98 VDD LPPFET W=0.62U L=0.12U M=1 
X2 VDD c hnet28 VDD LPPFET W=0.86U L=0.12U M=1 
X20 nmsi net86 nmin VDD LPPFET W=1.22U L=0.12U M=1 
X21 net128 cn m VDD LPPFET W=2.62U L=0.12U M=1 
X22 cn CK VSS VSS LPNFET W=0.48U L=0.12U M=1 
X23 nmsi net135 nmin VSS LPNFET W=0.88U L=0.12U M=1 
X24 net128 c m VSS LPNFET W=1.5U L=0.12U M=1 
X25 hnet46 s VSS VSS LPNFET W=0.36U L=0.12U M=1 
X26 nmsi nmen hnet46 VSS LPNFET W=0.36U L=0.12U M=1 
X27 hnet48 net137 nmsi VDD LPPFET W=0.5U L=0.12U M=1 
X28 VDD s hnet48 VDD LPPFET W=0.5U L=0.12U M=1 
X29 hnet52 SI VSS VSS LPNFET W=0.22U L=0.12U M=1 
X3 hnet28 nmsi pm VDD LPPFET W=0.86U L=0.12U M=1 
X30 nmsi SE hnet52 VSS LPNFET W=0.22U L=0.12U M=1 
X31 hnet54 nmse nmsi VDD LPPFET W=0.3U L=0.12U M=1 
X32 VDD SI hnet54 VDD LPPFET W=0.3U L=0.12U M=1 
X33 hnet58 m VSS VSS LPNFET W=0.18U L=0.12U M=1 
X34 pm c hnet58 VSS LPNFET W=0.18U L=0.12U M=1 
X35 hnet60 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X36 VDD m hnet60 VDD LPPFET W=0.28U L=0.12U M=1 
X37 hnet64 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X38 net128 cn hnet64 VSS LPNFET W=0.2U L=0.12U M=1 
X39 hnet66 c net128 VDD LPPFET W=0.28U L=0.12U M=1 
X4 hnet36 cn VSS VSS LPNFET W=0.66U L=0.12U M=1 
X40 VDD s hnet66 VDD LPPFET W=0.28U L=0.12U M=1 
X41 VDD D nmin VDD LPPFET W=1.22U L=0.12U M=1 
X42 nmin D VSS VSS LPNFET W=0.88U L=0.12U M=1 
X43 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X44 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X45 VDD net86 net135 VDD LPPFET W=0.28U L=0.12U M=1 
X46 net135 net86 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X47 VDD nmen net137 VDD LPPFET W=0.28U L=0.12U M=1 
X48 net137 nmen VSS VSS LPNFET W=0.2U L=0.12U M=1 
X49 VDD pm m VDD LPPFET W=2.78U L=0.12U M=1 
X5 pm nmsi hnet36 VSS LPNFET W=0.66U L=0.12U M=1 
X50 m pm VSS VSS LPNFET W=1.56U L=0.12U M=1 
X51 VDD net128 s VDD LPPFET W=0.28U L=0.12U M=1 
X52 s net128 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X53 VDD net128 Q VDD LPPFET W=2.6U L=0.12U M=1 
X54 Q net128 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X55 VDD net147 c VDD LPPFET W=2.02U L=0.12U M=1 
X56 c net147 VSS VSS LPNFET W=0.72U L=0.12U M=1 
X57 VDD CK net147 VDD LPPFET W=0.54U L=0.12U M=1 
X58 net147 CK VSS VSS LPNFET W=0.54U L=0.12U M=1 
X6 hnet32 cn VSS VSS LPNFET W=0.66U L=0.12U M=1 
X7 pm nmsi hnet32 VSS LPNFET W=0.66U L=0.12U M=1 
X8 nmen SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X9 nmen E VSS VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS SEDFFHQX4TS 

**** 
*.SUBCKT SEDFFHQX8TS Q CK D E SE SI 
.SUBCKT SEDFFHQX8TS Q CK D E SE SI VSS VDD
X0 VDD c hnet31 VDD LPPFET W=0.86U L=0.12U M=1 
X1 hnet31 nmsi pm VDD LPPFET W=0.86U L=0.12U M=1 
X10 VDD SE hnet38 VDD LPPFET W=0.4U L=0.12U M=1 
X11 hnet38 E nmen VDD LPPFET W=0.4U L=0.12U M=1 
X12 hnet44 nmse VSS VSS LPNFET W=0.2U L=0.12U M=1 
X13 net86 E hnet44 VSS LPNFET W=0.2U L=0.12U M=1 
X14 VDD nmse net86 VDD LPPFET W=0.28U L=0.12U M=1 
X15 VDD E net86 VDD LPPFET W=0.28U L=0.12U M=1 
X16 cn c net89 VDD LPPFET W=0.62U L=0.12U M=1 
X17 net89 CK VDD VDD LPPFET W=0.84U L=0.12U M=1 
X18 net98 CK VDD VDD LPPFET W=0.72U L=0.12U M=1 
X19 cn c net98 VDD LPPFET W=0.62U L=0.12U M=1 
X2 VDD c hnet28 VDD LPPFET W=0.86U L=0.12U M=1 
X20 nmsi net86 nmin VDD LPPFET W=1.22U L=0.12U M=1 
X21 net128 cn m VDD LPPFET W=2.62U L=0.12U M=1 
X22 cn CK VSS VSS LPNFET W=0.48U L=0.12U M=1 
X23 nmsi net135 nmin VSS LPNFET W=0.88U L=0.12U M=1 
X24 net128 c m VSS LPNFET W=1.5U L=0.12U M=1 
X25 hnet46 s VSS VSS LPNFET W=0.36U L=0.12U M=1 
X26 nmsi nmen hnet46 VSS LPNFET W=0.36U L=0.12U M=1 
X27 hnet48 net137 nmsi VDD LPPFET W=0.5U L=0.12U M=1 
X28 VDD s hnet48 VDD LPPFET W=0.5U L=0.12U M=1 
X29 hnet52 SI VSS VSS LPNFET W=0.22U L=0.12U M=1 
X3 hnet28 nmsi pm VDD LPPFET W=0.86U L=0.12U M=1 
X30 nmsi SE hnet52 VSS LPNFET W=0.22U L=0.12U M=1 
X31 hnet54 nmse nmsi VDD LPPFET W=0.3U L=0.12U M=1 
X32 VDD SI hnet54 VDD LPPFET W=0.3U L=0.12U M=1 
X33 hnet58 m VSS VSS LPNFET W=0.18U L=0.12U M=1 
X34 pm c hnet58 VSS LPNFET W=0.18U L=0.12U M=1 
X35 hnet60 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X36 VDD m hnet60 VDD LPPFET W=0.28U L=0.12U M=1 
X37 hnet64 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X38 net128 cn hnet64 VSS LPNFET W=0.2U L=0.12U M=1 
X39 hnet66 c net128 VDD LPPFET W=0.28U L=0.12U M=1 
X4 hnet36 cn VSS VSS LPNFET W=0.66U L=0.12U M=1 
X40 VDD s hnet66 VDD LPPFET W=0.28U L=0.12U M=1 
X41 VDD D nmin VDD LPPFET W=1.22U L=0.12U M=1 
X42 nmin D VSS VSS LPNFET W=0.88U L=0.12U M=1 
X43 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X44 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X45 VDD net86 net135 VDD LPPFET W=0.28U L=0.12U M=1 
X46 net135 net86 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X47 VDD nmen net137 VDD LPPFET W=0.28U L=0.12U M=1 
X48 net137 nmen VSS VSS LPNFET W=0.2U L=0.12U M=1 
X49 VDD pm m VDD LPPFET W=2.78U L=0.12U M=1 
X5 pm nmsi hnet36 VSS LPNFET W=0.66U L=0.12U M=1 
X50 m pm VSS VSS LPNFET W=1.56U L=0.12U M=1 
X51 VDD net128 s VDD LPPFET W=0.28U L=0.12U M=1 
X52 s net128 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X53 VDD net128 Q VDD LPPFET W=5.2U L=0.12U M=1 
X54 Q net128 VSS VSS LPNFET W=3.68U L=0.12U M=1 
X55 VDD net147 c VDD LPPFET W=2.02U L=0.12U M=1 
X56 c net147 VSS VSS LPNFET W=0.72U L=0.12U M=1 
X57 VDD CK net147 VDD LPPFET W=0.54U L=0.12U M=1 
X58 net147 CK VSS VSS LPNFET W=0.54U L=0.12U M=1 
X6 hnet32 cn VSS VSS LPNFET W=0.66U L=0.12U M=1 
X7 pm nmsi hnet32 VSS LPNFET W=0.66U L=0.12U M=1 
X8 nmen SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X9 nmen E VSS VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS SEDFFHQX8TS 

**** 
*.SUBCKT SEDFFTRX1TS Q QN CK D E RN SE SI 
.SUBCKT SEDFFTRX1TS Q QN CK D E RN SE SI VSS VDD
X0 nmrs SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X1 nmrs RN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X10 hnet46 c net130 VDD LPPFET W=0.26U L=0.12U M=1 
X11 VDD s hnet46 VDD LPPFET W=0.26U L=0.12U M=1 
X12 net103 net139 net112 VDD LPPFET W=0.36U L=0.12U M=1 
X13 net130 cn net153 VDD LPPFET W=0.64U L=0.12U M=1 
X14 net103 nmrs VDD VDD LPPFET W=0.36U L=0.12U M=1 
X15 net112 c pm VDD LPPFET W=0.36U L=0.12U M=1 
X16 net139 nmse nmsi VDD LPPFET W=0.28U L=0.12U M=1 
X17 net139 net167 net145 VDD LPPFET W=0.4U L=0.12U M=1 
X18 net145 net171 s VDD LPPFET W=0.44U L=0.12U M=1 
X19 net145 nmen nmin VDD LPPFET W=0.44U L=0.12U M=1 
X2 VDD SE hnet34 VDD LPPFET W=0.36U L=0.12U M=1 
X20 net127 nmrs VSS VSS LPNFET W=0.38U L=0.12U M=1 
X21 net130 c net153 VSS LPNFET W=0.46U L=0.12U M=1 
X22 net127 net139 VSS VSS LPNFET W=0.26U L=0.12U M=1 
X23 pm cn net127 VSS LPNFET W=0.26U L=0.12U M=1 
X24 net139 net167 nmsi VSS LPNFET W=0.2U L=0.12U M=1 
X25 net139 nmse net145 VSS LPNFET W=0.32U L=0.12U M=1 
X26 net145 nmen s VSS LPNFET W=0.32U L=0.12U M=1 
X27 net145 net171 nmin VSS LPNFET W=0.32U L=0.12U M=1 
X28 VDD s net149 VDD LPPFET W=0.28U L=0.12U M=1 
X29 net149 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 hnet34 RN nmrs VDD LPPFET W=0.36U L=0.12U M=1 
X30 VDD net149 QN VDD LPPFET W=0.64U L=0.12U M=1 
X31 QN net149 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X32 VDD m net153 VDD LPPFET W=0.64U L=0.12U M=1 
X33 net153 m VSS VSS LPNFET W=0.46U L=0.12U M=1 
X34 VDD pm m VDD LPPFET W=0.28U L=0.12U M=1 
X35 m pm VSS VSS LPNFET W=0.2U L=0.12U M=1 
X36 VDD net130 s VDD LPPFET W=0.8U L=0.12U M=1 
X37 s net130 VSS VSS LPNFET W=0.58U L=0.12U M=1 
X38 VDD s Q VDD LPPFET W=0.64U L=0.12U M=1 
X39 Q s VSS VSS LPNFET W=0.46U L=0.12U M=1 
X4 hnet38 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X40 VDD cn c VDD LPPFET W=0.3U L=0.12U M=1 
X41 c cn VSS VSS LPNFET W=0.22U L=0.12U M=1 
X42 VDD CK cn VDD LPPFET W=0.44U L=0.12U M=1 
X43 cn CK VSS VSS LPNFET W=0.32U L=0.12U M=1 
X44 VDD SI nmsi VDD LPPFET W=0.28U L=0.12U M=1 
X45 nmsi SI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X46 VDD nmse net167 VDD LPPFET W=0.28U L=0.12U M=1 
X47 net167 nmse VSS VSS LPNFET W=0.2U L=0.12U M=1 
X48 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X49 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X5 pm c hnet38 VSS LPNFET W=0.2U L=0.12U M=1 
X50 VDD nmen net171 VDD LPPFET W=0.28U L=0.12U M=1 
X51 net171 nmen VSS VSS LPNFET W=0.2U L=0.12U M=1 
X52 VDD E nmen VDD LPPFET W=0.28U L=0.12U M=1 
X53 nmen E VSS VSS LPNFET W=0.2U L=0.12U M=1 
X54 VDD D nmin VDD LPPFET W=0.44U L=0.12U M=1 
X55 nmin D VSS VSS LPNFET W=0.32U L=0.12U M=1 
X6 hnet40 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X7 VDD m hnet40 VDD LPPFET W=0.28U L=0.12U M=1 
X8 hnet44 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X9 net130 cn hnet44 VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS SEDFFTRX1TS 

**** 
*.SUBCKT SEDFFTRX2TS Q QN CK D E RN SE SI 
.SUBCKT SEDFFTRX2TS Q QN CK D E RN SE SI VSS VDD
X0 nmrs SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X1 nmrs RN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X10 hnet46 c net130 VDD LPPFET W=0.26U L=0.12U M=1 
X11 VDD s hnet46 VDD LPPFET W=0.26U L=0.12U M=1 
X12 net103 net139 net112 VDD LPPFET W=0.36U L=0.12U M=1 
X13 net130 cn net153 VDD LPPFET W=0.84U L=0.12U M=1 
X14 net103 nmrs VDD VDD LPPFET W=0.36U L=0.12U M=1 
X15 net112 c pm VDD LPPFET W=0.36U L=0.12U M=1 
X16 net139 nmse nmsi VDD LPPFET W=0.28U L=0.12U M=1 
X17 net139 net167 net145 VDD LPPFET W=0.44U L=0.12U M=1 
X18 net145 net171 s VDD LPPFET W=0.44U L=0.12U M=1 
X19 net145 nmen nmin VDD LPPFET W=0.44U L=0.12U M=1 
X2 VDD SE hnet34 VDD LPPFET W=0.36U L=0.12U M=1 
X20 net127 nmrs VSS VSS LPNFET W=0.38U L=0.12U M=1 
X21 net130 c net153 VSS LPNFET W=0.6U L=0.12U M=1 
X22 net127 net139 VSS VSS LPNFET W=0.26U L=0.12U M=1 
X23 pm cn net127 VSS LPNFET W=0.26U L=0.12U M=1 
X24 net139 net167 nmsi VSS LPNFET W=0.2U L=0.12U M=1 
X25 net139 nmse net145 VSS LPNFET W=0.32U L=0.12U M=1 
X26 net145 nmen s VSS LPNFET W=0.32U L=0.12U M=1 
X27 net145 net171 nmin VSS LPNFET W=0.32U L=0.12U M=1 
X28 VDD s net149 VDD LPPFET W=0.3U L=0.12U M=1 
X29 net149 s VSS VSS LPNFET W=0.22U L=0.12U M=1 
X3 hnet34 RN nmrs VDD LPPFET W=0.36U L=0.12U M=1 
X30 VDD net149 QN VDD LPPFET W=1.28U L=0.12U M=1 
X31 QN net149 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X32 VDD m net153 VDD LPPFET W=0.84U L=0.12U M=1 
X33 net153 m VSS VSS LPNFET W=0.56U L=0.12U M=1 
X34 VDD pm m VDD LPPFET W=0.28U L=0.12U M=1 
X35 m pm VSS VSS LPNFET W=0.24U L=0.12U M=1 
X36 VDD net130 s VDD LPPFET W=0.98U L=0.12U M=1 
X37 s net130 VSS VSS LPNFET W=0.7U L=0.12U M=1 
X38 VDD s Q VDD LPPFET W=1.28U L=0.12U M=1 
X39 Q s VSS VSS LPNFET W=0.92U L=0.12U M=1 
X4 hnet38 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X40 VDD cn c VDD LPPFET W=0.34U L=0.12U M=1 
X41 c cn VSS VSS LPNFET W=0.24U L=0.12U M=1 
X42 VDD CK cn VDD LPPFET W=0.5U L=0.12U M=1 
X43 cn CK VSS VSS LPNFET W=0.36U L=0.12U M=1 
X44 VDD SI nmsi VDD LPPFET W=0.28U L=0.12U M=1 
X45 nmsi SI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X46 VDD nmse net167 VDD LPPFET W=0.28U L=0.12U M=1 
X47 net167 nmse VSS VSS LPNFET W=0.2U L=0.12U M=1 
X48 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X49 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X5 pm c hnet38 VSS LPNFET W=0.2U L=0.12U M=1 
X50 VDD nmen net171 VDD LPPFET W=0.28U L=0.12U M=1 
X51 net171 nmen VSS VSS LPNFET W=0.2U L=0.12U M=1 
X52 VDD E nmen VDD LPPFET W=0.28U L=0.12U M=1 
X53 nmen E VSS VSS LPNFET W=0.2U L=0.12U M=1 
X54 VDD D nmin VDD LPPFET W=0.44U L=0.12U M=1 
X55 nmin D VSS VSS LPNFET W=0.32U L=0.12U M=1 
X6 hnet40 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X7 VDD m hnet40 VDD LPPFET W=0.28U L=0.12U M=1 
X8 hnet44 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X9 net130 cn hnet44 VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS SEDFFTRX2TS 

**** 
*.SUBCKT SEDFFTRX4TS Q QN CK D E RN SE SI 
.SUBCKT SEDFFTRX4TS Q QN CK D E RN SE SI VSS VDD
X0 nmrs SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X1 nmrs RN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X10 hnet46 c net130 VDD LPPFET W=0.26U L=0.12U M=1 
X11 VDD s hnet46 VDD LPPFET W=0.26U L=0.12U M=1 
X12 net103 net139 net112 VDD LPPFET W=0.36U L=0.12U M=1 
X13 net130 cn net153 VDD LPPFET W=1.2U L=0.12U M=1 
X14 net103 nmrs VDD VDD LPPFET W=0.36U L=0.12U M=1 
X15 net112 c pm VDD LPPFET W=0.36U L=0.12U M=1 
X16 net139 nmse nmsi VDD LPPFET W=0.28U L=0.12U M=1 
X17 net139 net167 net145 VDD LPPFET W=0.44U L=0.12U M=1 
X18 net145 net171 s VDD LPPFET W=0.44U L=0.12U M=1 
X19 net145 nmen nmin VDD LPPFET W=0.44U L=0.12U M=1 
X2 VDD SE hnet34 VDD LPPFET W=0.36U L=0.12U M=1 
X20 net127 nmrs VSS VSS LPNFET W=0.38U L=0.12U M=1 
X21 net130 c net153 VSS LPNFET W=0.9U L=0.12U M=1 
X22 net127 net139 VSS VSS LPNFET W=0.26U L=0.12U M=1 
X23 pm cn net127 VSS LPNFET W=0.26U L=0.12U M=1 
X24 net139 net167 nmsi VSS LPNFET W=0.2U L=0.12U M=1 
X25 net139 nmse net145 VSS LPNFET W=0.32U L=0.12U M=1 
X26 net145 nmen s VSS LPNFET W=0.32U L=0.12U M=1 
X27 net145 net171 nmin VSS LPNFET W=0.32U L=0.12U M=1 
X28 VDD s net149 VDD LPPFET W=0.62U L=0.12U M=1 
X29 net149 s VSS VSS LPNFET W=0.44U L=0.12U M=1 
X3 hnet34 RN nmrs VDD LPPFET W=0.36U L=0.12U M=1 
X30 VDD net149 QN VDD LPPFET W=2.56U L=0.12U M=1 
X31 QN net149 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X32 VDD m net153 VDD LPPFET W=1.2U L=0.12U M=1 
X33 net153 m VSS VSS LPNFET W=0.6U L=0.12U M=1 
X34 VDD pm m VDD LPPFET W=0.44U L=0.12U M=1 
X35 m pm VSS VSS LPNFET W=0.32U L=0.12U M=1 
X36 VDD net130 s VDD LPPFET W=1.56U L=0.12U M=1 
X37 s net130 VSS VSS LPNFET W=1.12U L=0.12U M=1 
X38 VDD s Q VDD LPPFET W=2.56U L=0.12U M=1 
X39 Q s VSS VSS LPNFET W=1.84U L=0.12U M=1 
X4 hnet38 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X40 VDD cn c VDD LPPFET W=0.42U L=0.12U M=1 
X41 c cn VSS VSS LPNFET W=0.3U L=0.12U M=1 
X42 VDD CK cn VDD LPPFET W=0.64U L=0.12U M=1 
X43 cn CK VSS VSS LPNFET W=0.42U L=0.12U M=1 
X44 VDD SI nmsi VDD LPPFET W=0.28U L=0.12U M=1 
X45 nmsi SI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X46 VDD nmse net167 VDD LPPFET W=0.28U L=0.12U M=1 
X47 net167 nmse VSS VSS LPNFET W=0.2U L=0.12U M=1 
X48 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X49 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X5 pm c hnet38 VSS LPNFET W=0.2U L=0.12U M=1 
X50 VDD nmen net171 VDD LPPFET W=0.28U L=0.12U M=1 
X51 net171 nmen VSS VSS LPNFET W=0.2U L=0.12U M=1 
X52 VDD E nmen VDD LPPFET W=0.28U L=0.12U M=1 
X53 nmen E VSS VSS LPNFET W=0.2U L=0.12U M=1 
X54 VDD D nmin VDD LPPFET W=0.44U L=0.12U M=1 
X55 nmin D VSS VSS LPNFET W=0.32U L=0.12U M=1 
X6 hnet40 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X7 VDD m hnet40 VDD LPPFET W=0.28U L=0.12U M=1 
X8 hnet44 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X9 net130 cn hnet44 VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS SEDFFTRX4TS 

**** 
*.SUBCKT SEDFFTRXLTS Q QN CK D E RN SE SI 
.SUBCKT SEDFFTRXLTS Q QN CK D E RN SE SI VSS VDD
X0 nmrs SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X1 nmrs RN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X10 hnet46 c net130 VDD LPPFET W=0.28U L=0.12U M=1 
X11 VDD s hnet46 VDD LPPFET W=0.28U L=0.12U M=1 
X12 net103 net139 net112 VDD LPPFET W=0.36U L=0.12U M=1 
X13 net130 cn net153 VDD LPPFET W=0.52U L=0.12U M=1 
X14 net103 nmrs VDD VDD LPPFET W=0.36U L=0.12U M=1 
X15 net112 c pm VDD LPPFET W=0.36U L=0.12U M=1 
X16 net139 nmse nmsi VDD LPPFET W=0.28U L=0.12U M=1 
X17 net139 net167 net145 VDD LPPFET W=0.4U L=0.12U M=1 
X18 net145 net171 s VDD LPPFET W=0.44U L=0.12U M=1 
X19 net145 nmen nmin VDD LPPFET W=0.44U L=0.12U M=1 
X2 VDD SE hnet34 VDD LPPFET W=0.36U L=0.12U M=1 
X20 net127 nmrs VSS VSS LPNFET W=0.38U L=0.12U M=1 
X21 net130 c net153 VSS LPNFET W=0.38U L=0.12U M=1 
X22 net127 net139 VSS VSS LPNFET W=0.26U L=0.12U M=1 
X23 pm cn net127 VSS LPNFET W=0.26U L=0.12U M=1 
X24 net139 net167 nmsi VSS LPNFET W=0.2U L=0.12U M=1 
X25 net139 nmse net145 VSS LPNFET W=0.32U L=0.12U M=1 
X26 net145 nmen s VSS LPNFET W=0.32U L=0.12U M=1 
X27 net145 net171 nmin VSS LPNFET W=0.32U L=0.12U M=1 
X28 VDD s net149 VDD LPPFET W=0.28U L=0.12U M=1 
X29 net149 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 hnet34 RN nmrs VDD LPPFET W=0.36U L=0.12U M=1 
X30 VDD net149 QN VDD LPPFET W=0.34U L=0.12U M=1 
X31 QN net149 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X32 VDD m net153 VDD LPPFET W=0.52U L=0.12U M=1 
X33 net153 m VSS VSS LPNFET W=0.38U L=0.12U M=1 
X34 VDD pm m VDD LPPFET W=0.28U L=0.12U M=1 
X35 m pm VSS VSS LPNFET W=0.2U L=0.12U M=1 
X36 VDD net130 s VDD LPPFET W=0.66U L=0.12U M=1 
X37 s net130 VSS VSS LPNFET W=0.48U L=0.12U M=1 
X38 VDD s Q VDD LPPFET W=0.34U L=0.12U M=1 
X39 Q s VSS VSS LPNFET W=0.24U L=0.12U M=1 
X4 hnet38 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X40 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X41 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X42 VDD CK cn VDD LPPFET W=0.44U L=0.12U M=1 
X43 cn CK VSS VSS LPNFET W=0.3U L=0.12U M=1 
X44 VDD SI nmsi VDD LPPFET W=0.28U L=0.12U M=1 
X45 nmsi SI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X46 VDD nmse net167 VDD LPPFET W=0.28U L=0.12U M=1 
X47 net167 nmse VSS VSS LPNFET W=0.2U L=0.12U M=1 
X48 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X49 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X5 pm c hnet38 VSS LPNFET W=0.2U L=0.12U M=1 
X50 VDD nmen net171 VDD LPPFET W=0.28U L=0.12U M=1 
X51 net171 nmen VSS VSS LPNFET W=0.2U L=0.12U M=1 
X52 VDD E nmen VDD LPPFET W=0.28U L=0.12U M=1 
X53 nmen E VSS VSS LPNFET W=0.2U L=0.12U M=1 
X54 VDD D nmin VDD LPPFET W=0.44U L=0.12U M=1 
X55 nmin D VSS VSS LPNFET W=0.32U L=0.12U M=1 
X6 hnet40 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X7 VDD m hnet40 VDD LPPFET W=0.28U L=0.12U M=1 
X8 hnet44 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X9 net130 cn hnet44 VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS SEDFFTRXLTS 

**** 
*.SUBCKT SEDFFX1TS Q QN CK D E SE SI 
.SUBCKT SEDFFX1TS Q QN CK D E SE SI VSS VDD
X0 hnet31 SI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X1 net71 SE hnet31 VSS LPNFET W=0.2U L=0.12U M=1 
X10 net102 SE VDD VDD LPPFET W=0.28U L=0.12U M=1 
X11 net108 E net102 VDD LPPFET W=0.28U L=0.12U M=1 
X12 net105 nmen net102 VDD LPPFET W=0.28U L=0.12U M=1 
X13 net74 D net105 VDD LPPFET W=0.28U L=0.12U M=1 
X14 net74 s net108 VDD LPPFET W=0.28U L=0.12U M=1 
X15 pm c net74 VDD LPPFET W=0.28U L=0.12U M=1 
X16 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X17 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X18 VDD E nmen VDD LPPFET W=0.28U L=0.12U M=1 
X19 nmen E VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 VDD SI hnet35 VDD LPPFET W=0.28U L=0.12U M=1 
X20 VDD net130 Q VDD LPPFET W=0.64U L=0.12U M=1 
X21 Q net130 VSS VSS LPNFET W=0.44U L=0.12U M=1 
X22 VDD s QN VDD LPPFET W=0.64U L=0.12U M=1 
X23 QN s VSS VSS LPNFET W=0.46U L=0.12U M=1 
X24 VDD net130 s VDD LPPFET W=0.28U L=0.12U M=1 
X25 s net130 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X26 VDD pm m VDD LPPFET W=0.28U L=0.12U M=1 
X27 m pm VSS VSS LPNFET W=0.2U L=0.12U M=1 
X28 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X29 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 hnet35 nmse net74 VDD LPPFET W=0.28U L=0.12U M=1 
X30 VDD CK cn VDD LPPFET W=0.3U L=0.12U M=1 
X31 cn CK VSS VSS LPNFET W=0.22U L=0.12U M=1 
X32 hnet53 m VSS VSS LPNFET W=0.22U L=0.12U M=1 
X33 net130 c hnet53 VSS LPNFET W=0.22U L=0.12U M=1 
X34 hnet55 cn net130 VDD LPPFET W=0.3U L=0.12U M=1 
X35 VDD m hnet55 VDD LPPFET W=0.3U L=0.12U M=1 
X36 hnet59 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X37 net130 cn hnet59 VSS LPNFET W=0.2U L=0.12U M=1 
X38 hnet61 c net130 VDD LPPFET W=0.28U L=0.12U M=1 
X39 VDD s hnet61 VDD LPPFET W=0.28U L=0.12U M=1 
X4 net79 nmse VSS VSS LPNFET W=0.2U L=0.12U M=1 
X40 hnet65 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X41 pm c hnet65 VSS LPNFET W=0.2U L=0.12U M=1 
X42 hnet67 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X43 VDD m hnet67 VDD LPPFET W=0.28U L=0.12U M=1 
X5 net82 nmen net79 VSS LPNFET W=0.2U L=0.12U M=1 
X6 net71 s net82 VSS LPNFET W=0.2U L=0.12U M=1 
X7 net88 E net79 VSS LPNFET W=0.2U L=0.12U M=1 
X8 net71 D net88 VSS LPNFET W=0.2U L=0.12U M=1 
X9 pm cn net71 VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS SEDFFX1TS 

**** 
*.SUBCKT SEDFFX2TS Q QN CK D E SE SI 
.SUBCKT SEDFFX2TS Q QN CK D E SE SI VSS VDD
X0 hnet31 SI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X1 net71 SE hnet31 VSS LPNFET W=0.2U L=0.12U M=1 
X10 net102 SE VDD VDD LPPFET W=0.28U L=0.12U M=1 
X11 net108 E net102 VDD LPPFET W=0.28U L=0.12U M=1 
X12 net105 nmen net102 VDD LPPFET W=0.28U L=0.12U M=1 
X13 net74 D net105 VDD LPPFET W=0.28U L=0.12U M=1 
X14 net74 s net108 VDD LPPFET W=0.28U L=0.12U M=1 
X15 pm c net74 VDD LPPFET W=0.28U L=0.12U M=1 
X16 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X17 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X18 VDD E nmen VDD LPPFET W=0.28U L=0.12U M=1 
X19 nmen E VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 VDD SI hnet35 VDD LPPFET W=0.28U L=0.12U M=1 
X20 VDD net130 Q VDD LPPFET W=1.28U L=0.12U M=1 
X21 Q net130 VSS VSS LPNFET W=0.88U L=0.12U M=1 
X22 VDD s QN VDD LPPFET W=1.26U L=0.12U M=1 
X23 QN s VSS VSS LPNFET W=0.9U L=0.12U M=1 
X24 VDD net130 s VDD LPPFET W=0.28U L=0.12U M=1 
X25 s net130 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X26 VDD pm m VDD LPPFET W=0.28U L=0.12U M=1 
X27 m pm VSS VSS LPNFET W=0.2U L=0.12U M=1 
X28 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X29 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 hnet35 nmse net74 VDD LPPFET W=0.28U L=0.12U M=1 
X30 VDD CK cn VDD LPPFET W=0.36U L=0.12U M=1 
X31 cn CK VSS VSS LPNFET W=0.26U L=0.12U M=1 
X32 hnet53 m VSS VSS LPNFET W=0.38U L=0.12U M=1 
X33 net130 c hnet53 VSS LPNFET W=0.38U L=0.12U M=1 
X34 hnet55 cn net130 VDD LPPFET W=0.52U L=0.12U M=1 
X35 VDD m hnet55 VDD LPPFET W=0.52U L=0.12U M=1 
X36 hnet59 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X37 net130 cn hnet59 VSS LPNFET W=0.2U L=0.12U M=1 
X38 hnet61 c net130 VDD LPPFET W=0.28U L=0.12U M=1 
X39 VDD s hnet61 VDD LPPFET W=0.28U L=0.12U M=1 
X4 net79 nmse VSS VSS LPNFET W=0.2U L=0.12U M=1 
X40 hnet65 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X41 pm c hnet65 VSS LPNFET W=0.2U L=0.12U M=1 
X42 hnet67 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X43 VDD m hnet67 VDD LPPFET W=0.28U L=0.12U M=1 
X5 net82 nmen net79 VSS LPNFET W=0.2U L=0.12U M=1 
X6 net71 s net82 VSS LPNFET W=0.2U L=0.12U M=1 
X7 net88 E net79 VSS LPNFET W=0.2U L=0.12U M=1 
X8 net71 D net88 VSS LPNFET W=0.2U L=0.12U M=1 
X9 pm cn net71 VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS SEDFFX2TS 

**** 
*.SUBCKT SEDFFX4TS Q QN CK D E SE SI 
.SUBCKT SEDFFX4TS Q QN CK D E SE SI VSS VDD
X0 hnet31 SI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X1 net71 SE hnet31 VSS LPNFET W=0.2U L=0.12U M=1 
X10 net102 SE VDD VDD LPPFET W=0.28U L=0.12U M=1 
X11 net108 E net102 VDD LPPFET W=0.28U L=0.12U M=1 
X12 net105 nmen net102 VDD LPPFET W=0.28U L=0.12U M=1 
X13 net74 D net105 VDD LPPFET W=0.28U L=0.12U M=1 
X14 net74 s net108 VDD LPPFET W=0.28U L=0.12U M=1 
X15 pm c net74 VDD LPPFET W=0.28U L=0.12U M=1 
X16 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X17 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X18 VDD E nmen VDD LPPFET W=0.28U L=0.12U M=1 
X19 nmen E VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 VDD SI hnet35 VDD LPPFET W=0.28U L=0.12U M=1 
X20 VDD net130 Q VDD LPPFET W=2.28U L=0.12U M=1 
X21 Q net130 VSS VSS LPNFET W=1.36U L=0.12U M=1 
X22 VDD s QN VDD LPPFET W=2.52U L=0.12U M=1 
X23 QN s VSS VSS LPNFET W=1.8U L=0.12U M=1 
X24 VDD net130 s VDD LPPFET W=0.52U L=0.12U M=1 
X25 s net130 VSS VSS LPNFET W=0.32U L=0.12U M=1 
X26 VDD pm m VDD LPPFET W=0.28U L=0.12U M=1 
X27 m pm VSS VSS LPNFET W=0.2U L=0.12U M=1 
X28 VDD cn c VDD LPPFET W=0.34U L=0.12U M=1 
X29 c cn VSS VSS LPNFET W=0.24U L=0.12U M=1 
X3 hnet35 nmse net74 VDD LPPFET W=0.28U L=0.12U M=1 
X30 VDD CK cn VDD LPPFET W=0.48U L=0.12U M=1 
X31 cn CK VSS VSS LPNFET W=0.32U L=0.12U M=1 
X32 hnet53 m VSS VSS LPNFET W=0.7U L=0.12U M=1 
X33 net130 c hnet53 VSS LPNFET W=0.7U L=0.12U M=1 
X34 hnet55 cn net130 VDD LPPFET W=0.96U L=0.12U M=1 
X35 VDD m hnet55 VDD LPPFET W=0.96U L=0.12U M=1 
X36 hnet59 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X37 net130 cn hnet59 VSS LPNFET W=0.2U L=0.12U M=1 
X38 hnet61 c net130 VDD LPPFET W=0.28U L=0.12U M=1 
X39 VDD s hnet61 VDD LPPFET W=0.28U L=0.12U M=1 
X4 net79 nmse VSS VSS LPNFET W=0.2U L=0.12U M=1 
X40 hnet65 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X41 pm c hnet65 VSS LPNFET W=0.2U L=0.12U M=1 
X42 hnet67 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X43 VDD m hnet67 VDD LPPFET W=0.28U L=0.12U M=1 
X5 net82 nmen net79 VSS LPNFET W=0.2U L=0.12U M=1 
X6 net71 s net82 VSS LPNFET W=0.2U L=0.12U M=1 
X7 net88 E net79 VSS LPNFET W=0.2U L=0.12U M=1 
X8 net71 D net88 VSS LPNFET W=0.2U L=0.12U M=1 
X9 pm cn net71 VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS SEDFFX4TS 

**** 
*.SUBCKT SEDFFXLTS Q QN CK D E SE SI 
.SUBCKT SEDFFXLTS Q QN CK D E SE SI VSS VDD
X0 hnet31 SI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X1 net71 SE hnet31 VSS LPNFET W=0.2U L=0.12U M=1 
X10 net102 SE VDD VDD LPPFET W=0.28U L=0.12U M=1 
X11 net108 E net102 VDD LPPFET W=0.28U L=0.12U M=1 
X12 net105 nmen net102 VDD LPPFET W=0.28U L=0.12U M=1 
X13 net74 D net105 VDD LPPFET W=0.28U L=0.12U M=1 
X14 net74 s net108 VDD LPPFET W=0.28U L=0.12U M=1 
X15 pm c net74 VDD LPPFET W=0.28U L=0.12U M=1 
X16 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X17 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X18 VDD E nmen VDD LPPFET W=0.28U L=0.12U M=1 
X19 nmen E VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 VDD SI hnet35 VDD LPPFET W=0.28U L=0.12U M=1 
X20 VDD net130 Q VDD LPPFET W=0.34U L=0.12U M=1 
X21 Q net130 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X22 VDD s QN VDD LPPFET W=0.34U L=0.12U M=1 
X23 QN s VSS VSS LPNFET W=0.24U L=0.12U M=1 
X24 VDD net130 s VDD LPPFET W=0.28U L=0.12U M=1 
X25 s net130 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X26 VDD pm m VDD LPPFET W=0.28U L=0.12U M=1 
X27 m pm VSS VSS LPNFET W=0.2U L=0.12U M=1 
X28 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X29 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 hnet35 nmse net74 VDD LPPFET W=0.28U L=0.12U M=1 
X30 VDD CK cn VDD LPPFET W=0.3U L=0.12U M=1 
X31 cn CK VSS VSS LPNFET W=0.22U L=0.12U M=1 
X32 hnet53 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X33 net130 c hnet53 VSS LPNFET W=0.2U L=0.12U M=1 
X34 hnet55 cn net130 VDD LPPFET W=0.28U L=0.12U M=1 
X35 VDD m hnet55 VDD LPPFET W=0.28U L=0.12U M=1 
X36 hnet59 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X37 net130 cn hnet59 VSS LPNFET W=0.2U L=0.12U M=1 
X38 hnet61 c net130 VDD LPPFET W=0.28U L=0.12U M=1 
X39 VDD s hnet61 VDD LPPFET W=0.28U L=0.12U M=1 
X4 net79 nmse VSS VSS LPNFET W=0.2U L=0.12U M=1 
X40 hnet65 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X41 pm c hnet65 VSS LPNFET W=0.2U L=0.12U M=1 
X42 hnet67 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X43 VDD m hnet67 VDD LPPFET W=0.28U L=0.12U M=1 
X5 net82 nmen net79 VSS LPNFET W=0.2U L=0.12U M=1 
X6 net71 s net82 VSS LPNFET W=0.2U L=0.12U M=1 
X7 net88 E net79 VSS LPNFET W=0.2U L=0.12U M=1 
X8 net71 D net88 VSS LPNFET W=0.2U L=0.12U M=1 
X9 pm cn net71 VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS SEDFFXLTS 

**** 
*.SUBCKT SMDFFHQX1TS Q CK D0 D1 S0 SE SI 
.SUBCKT SMDFFHQX1TS Q CK D0 D1 S0 SE SI VSS VDD
X0 nmsel SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X1 nmsel S0 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X10 hnet43 cn VSS VSS LPNFET W=0.42U L=0.12U M=1 
X11 pm nmsi hnet43 VSS LPNFET W=0.42U L=0.12U M=1 
X12 net92 CK VDD VDD LPPFET W=0.7U L=0.12U M=1 
X13 cn c net92 VDD LPPFET W=0.52U L=0.12U M=1 
X14 nmsi net135 nmin0 VDD LPPFET W=0.38U L=0.12U M=1 
X15 nmsi net80 nmin1 VDD LPPFET W=0.38U L=0.12U M=1 
X16 net124 cn m VDD LPPFET W=0.96U L=0.12U M=1 
X17 cn CK VSS VSS LPNFET W=0.2U L=0.12U M=1 
X18 nmsi nmsel nmin0 VSS LPNFET W=0.28U L=0.12U M=1 
X19 nmsi net133 nmin1 VSS LPNFET W=0.28U L=0.12U M=1 
X2 VDD SE hnet29 VDD LPPFET W=0.38U L=0.12U M=1 
X20 net124 c m VSS LPNFET W=0.5U L=0.12U M=1 
X21 hnet45 SI VSS VSS LPNFET W=0.2U L=0.12U M=1 
X22 nmsi SE hnet45 VSS LPNFET W=0.2U L=0.12U M=1 
X23 hnet47 nmse nmsi VDD LPPFET W=0.28U L=0.12U M=1 
X24 VDD SI hnet47 VDD LPPFET W=0.28U L=0.12U M=1 
X25 hnet51 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X26 pm c hnet51 VSS LPNFET W=0.2U L=0.12U M=1 
X27 hnet53 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X28 VDD m hnet53 VDD LPPFET W=0.28U L=0.12U M=1 
X29 hnet57 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 hnet29 S0 nmsel VDD LPPFET W=0.38U L=0.12U M=1 
X30 net124 cn hnet57 VSS LPNFET W=0.2U L=0.12U M=1 
X31 hnet59 c net124 VDD LPPFET W=0.28U L=0.12U M=1 
X32 VDD s hnet59 VDD LPPFET W=0.28U L=0.12U M=1 
X33 VDD D0 nmin0 VDD LPPFET W=0.38U L=0.12U M=1 
X34 nmin0 D0 VSS VSS LPNFET W=0.28U L=0.12U M=1 
X35 VDD D1 nmin1 VDD LPPFET W=0.38U L=0.12U M=1 
X36 nmin1 D1 VSS VSS LPNFET W=0.28U L=0.12U M=1 
X37 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X38 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X39 VDD net80 net133 VDD LPPFET W=0.28U L=0.12U M=1 
X4 hnet35 nmse VSS VSS LPNFET W=0.2U L=0.12U M=1 
X40 net133 net80 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X41 VDD nmsel net135 VDD LPPFET W=0.28U L=0.12U M=1 
X42 net135 nmsel VSS VSS LPNFET W=0.2U L=0.12U M=1 
X43 VDD pm m VDD LPPFET W=0.96U L=0.12U M=1 
X44 m pm VSS VSS LPNFET W=0.5U L=0.12U M=1 
X45 VDD net124 s VDD LPPFET W=0.28U L=0.12U M=1 
X46 s net124 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X47 VDD net124 Q VDD LPPFET W=0.74U L=0.12U M=1 
X48 Q net124 VSS VSS LPNFET W=0.56U L=0.12U M=1 
X49 VDD net145 c VDD LPPFET W=0.84U L=0.12U M=1 
X5 net80 S0 hnet35 VSS LPNFET W=0.2U L=0.12U M=1 
X50 c net145 VSS VSS LPNFET W=0.3U L=0.12U M=1 
X51 VDD CK net145 VDD LPPFET W=0.28U L=0.12U M=1 
X52 net145 CK VSS VSS LPNFET W=0.28U L=0.12U M=1 
X6 VDD nmse net80 VDD LPPFET W=0.28U L=0.12U M=1 
X7 VDD S0 net80 VDD LPPFET W=0.28U L=0.12U M=1 
X8 VDD c hnet39 VDD LPPFET W=0.58U L=0.12U M=1 
X9 hnet39 nmsi pm VDD LPPFET W=0.58U L=0.12U M=1 
.ENDS SMDFFHQX1TS 

**** 
*.SUBCKT SMDFFHQX2TS Q CK D0 D1 S0 SE SI 
.SUBCKT SMDFFHQX2TS Q CK D0 D1 S0 SE SI VSS VDD
X0 nmsel SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X1 nmsel S0 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X10 hnet43 cn VSS VSS LPNFET W=0.66U L=0.12U M=1 
X11 pm nmsi hnet43 VSS LPNFET W=0.66U L=0.12U M=1 
X12 net92 CK VDD VDD LPPFET W=0.9U L=0.12U M=1 
X13 cn c net92 VDD LPPFET W=0.68U L=0.12U M=1 
X14 nmsi net135 nmin0 VDD LPPFET W=0.68U L=0.12U M=1 
X15 nmsi net80 nmin1 VDD LPPFET W=0.68U L=0.12U M=1 
X16 net124 cn m VDD LPPFET W=1.38U L=0.12U M=1 
X17 cn CK VSS VSS LPNFET W=0.28U L=0.12U M=1 
X18 nmsi nmsel nmin0 VSS LPNFET W=0.46U L=0.12U M=1 
X19 nmsi net133 nmin1 VSS LPNFET W=0.5U L=0.12U M=1 
X2 VDD SE hnet29 VDD LPPFET W=0.4U L=0.12U M=1 
X20 net124 c m VSS LPNFET W=0.7U L=0.12U M=1 
X21 hnet45 SI VSS VSS LPNFET W=0.24U L=0.12U M=1 
X22 nmsi SE hnet45 VSS LPNFET W=0.24U L=0.12U M=1 
X23 hnet47 nmse nmsi VDD LPPFET W=0.34U L=0.12U M=1 
X24 VDD SI hnet47 VDD LPPFET W=0.34U L=0.12U M=1 
X25 hnet51 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X26 pm c hnet51 VSS LPNFET W=0.2U L=0.12U M=1 
X27 hnet53 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X28 VDD m hnet53 VDD LPPFET W=0.28U L=0.12U M=1 
X29 hnet57 s VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 hnet29 S0 nmsel VDD LPPFET W=0.4U L=0.12U M=1 
X30 net124 cn hnet57 VSS LPNFET W=0.2U L=0.12U M=1 
X31 hnet59 c net124 VDD LPPFET W=0.28U L=0.12U M=1 
X32 VDD s hnet59 VDD LPPFET W=0.28U L=0.12U M=1 
X33 VDD D0 nmin0 VDD LPPFET W=0.68U L=0.12U M=1 
X34 nmin0 D0 VSS VSS LPNFET W=0.52U L=0.12U M=1 
X35 VDD D1 nmin1 VDD LPPFET W=0.68U L=0.12U M=1 
X36 nmin1 D1 VSS VSS LPNFET W=0.5U L=0.12U M=1 
X37 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X38 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X39 VDD net80 net133 VDD LPPFET W=0.28U L=0.12U M=1 
X4 hnet35 nmse VSS VSS LPNFET W=0.2U L=0.12U M=1 
X40 net133 net80 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X41 VDD nmsel net135 VDD LPPFET W=0.28U L=0.12U M=1 
X42 net135 nmsel VSS VSS LPNFET W=0.2U L=0.12U M=1 
X43 VDD pm m VDD LPPFET W=1.48U L=0.12U M=1 
X44 m pm VSS VSS LPNFET W=0.7U L=0.12U M=1 
X45 VDD net124 s VDD LPPFET W=0.28U L=0.12U M=1 
X46 s net124 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X47 VDD net124 Q VDD LPPFET W=1.48U L=0.12U M=1 
X48 Q net124 VSS VSS LPNFET W=0.72U L=0.12U M=1 
X49 VDD net145 c VDD LPPFET W=1.18U L=0.12U M=1 
X5 net80 S0 hnet35 VSS LPNFET W=0.2U L=0.12U M=1 
X50 c net145 VSS VSS LPNFET W=0.42U L=0.12U M=1 
X51 VDD CK net145 VDD LPPFET W=0.32U L=0.12U M=1 
X52 net145 CK VSS VSS LPNFET W=0.32U L=0.12U M=1 
X6 VDD nmse net80 VDD LPPFET W=0.28U L=0.12U M=1 
X7 VDD S0 net80 VDD LPPFET W=0.28U L=0.12U M=1 
X8 VDD c hnet39 VDD LPPFET W=1U L=0.12U M=1 
X9 hnet39 nmsi pm VDD LPPFET W=1U L=0.12U M=1 
.ENDS SMDFFHQX2TS 

**** 
*.SUBCKT SMDFFHQX4TS Q CK D0 D1 S0 SE SI 
.SUBCKT SMDFFHQX4TS Q CK D0 D1 S0 SE SI VSS VDD
X0 VDD c hnet33 VDD LPPFET W=0.9U L=0.12U M=1 
X1 hnet33 nmsi pm VDD LPPFET W=0.9U L=0.12U M=1 
X10 VDD SE hnet40 VDD LPPFET W=0.4U L=0.12U M=1 
X11 hnet40 S0 nmsel VDD LPPFET W=0.4U L=0.12U M=1 
X12 hnet46 nmse VSS VSS LPNFET W=0.24U L=0.12U M=1 
X13 net83 S0 hnet46 VSS LPNFET W=0.24U L=0.12U M=1 
X14 VDD nmse net83 VDD LPPFET W=0.28U L=0.12U M=1 
X15 VDD S0 net83 VDD LPPFET W=0.28U L=0.12U M=1 
X16 cn c net90 VDD LPPFET W=0.64U L=0.12U M=1 
X17 net90 CK VDD VDD LPPFET W=0.84U L=0.12U M=1 
X18 net93 CK VDD VDD LPPFET W=0.72U L=0.12U M=1 
X19 cn c net93 VDD LPPFET W=0.64U L=0.12U M=1 
X2 VDD c hnet30 VDD LPPFET W=0.9U L=0.12U M=1 
X20 nmsi net138 nmin0 VDD LPPFET W=1.22U L=0.12U M=1 
X21 nmsi net83 nmin1 VDD LPPFET W=1.22U L=0.12U M=1 
X22 net127 cn m VDD LPPFET W=2.72U L=0.12U M=1 
X23 cn CK VSS VSS LPNFET W=0.54U L=0.12U M=1 
X24 nmsi nmsel nmin0 VSS LPNFET W=0.88U L=0.12U M=1 
X25 nmsi net136 nmin1 VSS LPNFET W=0.88U L=0.12U M=1 
X26 net127 c m VSS LPNFET W=1.5U L=0.12U M=1 
X27 hnet48 SI VSS VSS LPNFET W=0.44U L=0.12U M=1 
X28 nmsi SE hnet48 VSS LPNFET W=0.44U L=0.12U M=1 
X29 hnet50 nmse nmsi VDD LPPFET W=0.62U L=0.12U M=1 
X3 hnet30 nmsi pm VDD LPPFET W=0.9U L=0.12U M=1 
X30 VDD SI hnet50 VDD LPPFET W=0.62U L=0.12U M=1 
X31 hnet54 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X32 pm c hnet54 VSS LPNFET W=0.2U L=0.12U M=1 
X33 hnet56 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X34 VDD m hnet56 VDD LPPFET W=0.28U L=0.12U M=1 
X35 hnet60 s VSS VSS LPNFET W=0.32U L=0.12U M=1 
X36 net127 cn hnet60 VSS LPNFET W=0.32U L=0.12U M=1 
X37 hnet62 c net127 VDD LPPFET W=0.28U L=0.12U M=1 
X38 VDD s hnet62 VDD LPPFET W=0.28U L=0.12U M=1 
X39 VDD D0 nmin0 VDD LPPFET W=1.22U L=0.12U M=1 
X4 hnet38 cn VSS VSS LPNFET W=0.66U L=0.12U M=1 
X40 nmin0 D0 VSS VSS LPNFET W=0.88U L=0.12U M=1 
X41 VDD D1 nmin1 VDD LPPFET W=1.22U L=0.12U M=1 
X42 nmin1 D1 VSS VSS LPNFET W=0.88U L=0.12U M=1 
X43 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X44 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X45 VDD net83 net136 VDD LPPFET W=0.28U L=0.12U M=1 
X46 net136 net83 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X47 VDD nmsel net138 VDD LPPFET W=0.28U L=0.12U M=1 
X48 net138 nmsel VSS VSS LPNFET W=0.2U L=0.12U M=1 
X49 VDD pm m VDD LPPFET W=2.72U L=0.12U M=1 
X5 pm nmsi hnet38 VSS LPNFET W=0.66U L=0.12U M=1 
X50 m pm VSS VSS LPNFET W=1.56U L=0.12U M=1 
X51 VDD net127 s VDD LPPFET W=0.28U L=0.12U M=1 
X52 s net127 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X53 VDD net127 Q VDD LPPFET W=2.6U L=0.12U M=1 
X54 Q net127 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X55 VDD net148 c VDD LPPFET W=2.02U L=0.12U M=1 
X56 c net148 VSS VSS LPNFET W=0.72U L=0.12U M=1 
X57 VDD CK net148 VDD LPPFET W=0.54U L=0.12U M=1 
X58 net148 CK VSS VSS LPNFET W=0.54U L=0.12U M=1 
X6 hnet34 cn VSS VSS LPNFET W=0.66U L=0.12U M=1 
X7 pm nmsi hnet34 VSS LPNFET W=0.66U L=0.12U M=1 
X8 nmsel SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X9 nmsel S0 VSS VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS SMDFFHQX4TS 

**** 
*.SUBCKT SMDFFHQX8TS Q CK D0 D1 S0 SE SI 
.SUBCKT SMDFFHQX8TS Q CK D0 D1 S0 SE SI VSS VDD
X0 VDD c hnet33 VDD LPPFET W=0.9U L=0.12U M=1 
X1 hnet33 nmsi pm VDD LPPFET W=0.9U L=0.12U M=1 
X10 VDD SE hnet40 VDD LPPFET W=0.4U L=0.12U M=1 
X11 hnet40 S0 nmsel VDD LPPFET W=0.4U L=0.12U M=1 
X12 hnet46 nmse VSS VSS LPNFET W=0.24U L=0.12U M=1 
X13 net83 S0 hnet46 VSS LPNFET W=0.24U L=0.12U M=1 
X14 VDD nmse net83 VDD LPPFET W=0.28U L=0.12U M=1 
X15 VDD S0 net83 VDD LPPFET W=0.28U L=0.12U M=1 
X16 cn c net90 VDD LPPFET W=0.64U L=0.12U M=1 
X17 net90 CK VDD VDD LPPFET W=0.84U L=0.12U M=1 
X18 net93 CK VDD VDD LPPFET W=0.72U L=0.12U M=1 
X19 cn c net93 VDD LPPFET W=0.64U L=0.12U M=1 
X2 VDD c hnet30 VDD LPPFET W=0.9U L=0.12U M=1 
X20 nmsi net138 nmin0 VDD LPPFET W=1.22U L=0.12U M=1 
X21 nmsi net83 nmin1 VDD LPPFET W=1.22U L=0.12U M=1 
X22 net127 cn m VDD LPPFET W=2.72U L=0.12U M=1 
X23 cn CK VSS VSS LPNFET W=0.54U L=0.12U M=1 
X24 nmsi nmsel nmin0 VSS LPNFET W=0.88U L=0.12U M=1 
X25 nmsi net136 nmin1 VSS LPNFET W=0.88U L=0.12U M=1 
X26 net127 c m VSS LPNFET W=1.5U L=0.12U M=1 
X27 hnet48 SI VSS VSS LPNFET W=0.44U L=0.12U M=1 
X28 nmsi SE hnet48 VSS LPNFET W=0.44U L=0.12U M=1 
X29 hnet50 nmse nmsi VDD LPPFET W=0.62U L=0.12U M=1 
X3 hnet30 nmsi pm VDD LPPFET W=0.9U L=0.12U M=1 
X30 VDD SI hnet50 VDD LPPFET W=0.62U L=0.12U M=1 
X31 hnet54 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X32 pm c hnet54 VSS LPNFET W=0.2U L=0.12U M=1 
X33 hnet56 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X34 VDD m hnet56 VDD LPPFET W=0.28U L=0.12U M=1 
X35 hnet60 s VSS VSS LPNFET W=0.32U L=0.12U M=1 
X36 net127 cn hnet60 VSS LPNFET W=0.32U L=0.12U M=1 
X37 hnet62 c net127 VDD LPPFET W=0.28U L=0.12U M=1 
X38 VDD s hnet62 VDD LPPFET W=0.28U L=0.12U M=1 
X39 VDD D0 nmin0 VDD LPPFET W=1.22U L=0.12U M=1 
X4 hnet38 cn VSS VSS LPNFET W=0.66U L=0.12U M=1 
X40 nmin0 D0 VSS VSS LPNFET W=0.88U L=0.12U M=1 
X41 VDD D1 nmin1 VDD LPPFET W=1.22U L=0.12U M=1 
X42 nmin1 D1 VSS VSS LPNFET W=0.88U L=0.12U M=1 
X43 VDD SE nmse VDD LPPFET W=0.28U L=0.12U M=1 
X44 nmse SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X45 VDD net83 net136 VDD LPPFET W=0.28U L=0.12U M=1 
X46 net136 net83 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X47 VDD nmsel net138 VDD LPPFET W=0.28U L=0.12U M=1 
X48 net138 nmsel VSS VSS LPNFET W=0.2U L=0.12U M=1 
X49 VDD pm m VDD LPPFET W=2.72U L=0.12U M=1 
X5 pm nmsi hnet38 VSS LPNFET W=0.66U L=0.12U M=1 
X50 m pm VSS VSS LPNFET W=1.56U L=0.12U M=1 
X51 VDD net127 s VDD LPPFET W=0.28U L=0.12U M=1 
X52 s net127 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X53 VDD net127 Q VDD LPPFET W=5.2U L=0.12U M=1 
X54 Q net127 VSS VSS LPNFET W=3.68U L=0.12U M=1 
X55 VDD net148 c VDD LPPFET W=2.02U L=0.12U M=1 
X56 c net148 VSS VSS LPNFET W=0.72U L=0.12U M=1 
X57 VDD CK net148 VDD LPPFET W=0.54U L=0.12U M=1 
X58 net148 CK VSS VSS LPNFET W=0.54U L=0.12U M=1 
X6 hnet34 cn VSS VSS LPNFET W=0.66U L=0.12U M=1 
X7 pm nmsi hnet34 VSS LPNFET W=0.66U L=0.12U M=1 
X8 nmsel SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X9 nmsel S0 VSS VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS SMDFFHQX8TS 

**** 
*.SUBCKT TBUFX12TS Y A OE 
.SUBCKT TBUFX12TS Y A OE VSS VDD
X0 VDD OE nmen VDD LPPFET W=0.52U L=0.12U M=1 
X1 nmen OE VSS VSS LPNFET W=0.38U L=0.12U M=1 
X2 net28 A VSS VSS LPNFET W=2.2U L=0.12U M=1 
X3 net28 nmen VSS VSS LPNFET W=0.64U L=0.12U M=1 
X4 Y net28 VSS VSS LPNFET W=5.52U L=0.12U M=1 
X5 nmin OE net28 VSS LPNFET W=1.14U L=0.12U M=1 
X6 nmin A VDD VDD LPPFET W=3.06U L=0.12U M=1 
X7 nmin OE VDD VDD LPPFET W=0.94U L=0.12U M=1 
X8 net28 nmen nmin VDD LPPFET W=1.54U L=0.12U M=1 
X9 Y nmin VDD VDD LPPFET W=7.32U L=0.12U M=1 
.ENDS TBUFX12TS 

**** 
*.SUBCKT TBUFX16TS Y A OE 
.SUBCKT TBUFX16TS Y A OE VSS VDD
X0 VDD OE nmen VDD LPPFET W=0.7U L=0.12U M=1 
X1 nmen OE VSS VSS LPNFET W=0.5U L=0.12U M=1 
X2 net28 A VSS VSS LPNFET W=2.7U L=0.12U M=1 
X3 net28 nmen VSS VSS LPNFET W=0.82U L=0.12U M=1 
X4 Y net28 VSS VSS LPNFET W=6.06U L=0.12U M=1 
X5 nmin OE net28 VSS LPNFET W=1.18U L=0.12U M=1 
X6 nmin A VDD VDD LPPFET W=3.9U L=0.12U M=1 
X7 nmin OE VDD VDD LPPFET W=1.26U L=0.12U M=1 
X8 net28 nmen nmin VDD LPPFET W=1.98U L=0.12U M=1 
X9 Y nmin VDD VDD LPPFET W=9.16U L=0.12U M=1 
.ENDS TBUFX16TS 

**** 
*.SUBCKT TBUFX1TS Y A OE 
.SUBCKT TBUFX1TS Y A OE VSS VDD
X0 VDD OE nmen VDD LPPFET W=0.28U L=0.12U M=1 
X1 nmen OE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 net28 A VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 net28 nmen VSS VSS LPNFET W=0.18U L=0.12U M=1 
X4 Y net28 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X5 nmin OE net28 VSS LPNFET W=0.2U L=0.12U M=1 
X6 nmin A VDD VDD LPPFET W=0.28U L=0.12U M=1 
X7 nmin OE VDD VDD LPPFET W=0.28U L=0.12U M=1 
X8 net28 nmen nmin VDD LPPFET W=0.28U L=0.12U M=1 
X9 Y nmin VDD VDD LPPFET W=0.64U L=0.12U M=1 
.ENDS TBUFX1TS 

**** 
*.SUBCKT TBUFX20TS Y A OE 
.SUBCKT TBUFX20TS Y A OE VSS VDD
X0 VDD OE nmen VDD LPPFET W=0.82U L=0.12U M=1 
X1 nmen OE VSS VSS LPNFET W=0.62U L=0.12U M=1 
X2 net28 A VSS VSS LPNFET W=3.24U L=0.12U M=1 
X3 net28 nmen VSS VSS LPNFET W=1.06U L=0.12U M=1 
X4 Y net28 VSS VSS LPNFET W=7.58U L=0.12U M=1 
X5 nmin OE net28 VSS LPNFET W=1.2U L=0.12U M=1 
X6 nmin A VDD VDD LPPFET W=4.44U L=0.12U M=1 
X7 nmin OE VDD VDD LPPFET W=1.6U L=0.12U M=1 
X8 net28 nmen nmin VDD LPPFET W=1.84U L=0.12U M=1 
X9 Y nmin VDD VDD LPPFET W=11.42U L=0.12U M=1 
.ENDS TBUFX20TS 

**** 
*.SUBCKT TBUFX2TS Y A OE 
.SUBCKT TBUFX2TS Y A OE VSS VDD
X0 VDD OE nmen VDD LPPFET W=0.28U L=0.12U M=1 
X1 nmen OE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 net28 A VSS VSS LPNFET W=0.36U L=0.12U M=1 
X3 net28 nmen VSS VSS LPNFET W=0.18U L=0.12U M=1 
X4 Y net28 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X5 nmin OE net28 VSS LPNFET W=0.2U L=0.12U M=1 
X6 nmin A VDD VDD LPPFET W=0.5U L=0.12U M=1 
X7 nmin OE VDD VDD LPPFET W=0.28U L=0.12U M=1 
X8 net28 nmen nmin VDD LPPFET W=0.28U L=0.12U M=1 
X9 Y nmin VDD VDD LPPFET W=1.24U L=0.12U M=1 
.ENDS TBUFX2TS 

**** 
*.SUBCKT TBUFX3TS Y A OE 
.SUBCKT TBUFX3TS Y A OE VSS VDD
X0 VDD OE nmen VDD LPPFET W=0.28U L=0.12U M=1 
X1 nmen OE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 net28 A VSS VSS LPNFET W=0.56U L=0.12U M=1 
X3 net28 nmen VSS VSS LPNFET W=0.18U L=0.12U M=1 
X4 Y net28 VSS VSS LPNFET W=1.32U L=0.12U M=1 
X5 nmin OE net28 VSS LPNFET W=0.28U L=0.12U M=1 
X6 nmin A VDD VDD LPPFET W=0.78U L=0.12U M=1 
X7 nmin OE VDD VDD LPPFET W=0.28U L=0.12U M=1 
X8 net28 nmen nmin VDD LPPFET W=0.38U L=0.12U M=1 
X9 Y nmin VDD VDD LPPFET W=1.92U L=0.12U M=1 
.ENDS TBUFX3TS 

**** 
*.SUBCKT TBUFX4TS Y A OE 
.SUBCKT TBUFX4TS Y A OE VSS VDD
X0 VDD OE nmen VDD LPPFET W=0.28U L=0.12U M=1 
X1 nmen OE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 net28 A VSS VSS LPNFET W=0.66U L=0.12U M=1 
X3 net28 nmen VSS VSS LPNFET W=0.22U L=0.12U M=1 
X4 Y net28 VSS VSS LPNFET W=1.76U L=0.12U M=1 
X5 nmin OE net28 VSS LPNFET W=0.36U L=0.12U M=1 
X6 nmin A VDD VDD LPPFET W=1.02U L=0.12U M=1 
X7 nmin OE VDD VDD LPPFET W=0.34U L=0.12U M=1 
X8 net28 nmen nmin VDD LPPFET W=0.5U L=0.12U M=1 
X9 Y nmin VDD VDD LPPFET W=2.56U L=0.12U M=1 
.ENDS TBUFX4TS 

**** 
*.SUBCKT TBUFX6TS Y A OE 
.SUBCKT TBUFX6TS Y A OE VSS VDD
X0 VDD OE nmen VDD LPPFET W=0.28U L=0.12U M=1 
X1 nmen OE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 net28 A VSS VSS LPNFET W=0.92U L=0.12U M=1 
X3 net28 nmen VSS VSS LPNFET W=0.34U L=0.12U M=1 
X4 Y net28 VSS VSS LPNFET W=2.7U L=0.12U M=1 
X5 nmin OE net28 VSS LPNFET W=0.56U L=0.12U M=1 
X6 nmin A VDD VDD LPPFET W=1.54U L=0.12U M=1 
X7 nmin OE VDD VDD LPPFET W=0.48U L=0.12U M=1 
X8 net28 nmen nmin VDD LPPFET W=0.78U L=0.12U M=1 
X9 Y nmin VDD VDD LPPFET W=3.5U L=0.12U M=1 
.ENDS TBUFX6TS 

**** 
*.SUBCKT TBUFX8TS Y A OE 
.SUBCKT TBUFX8TS Y A OE VSS VDD
X0 VDD OE nmen VDD LPPFET W=0.34U L=0.12U M=1 
X1 nmen OE VSS VSS LPNFET W=0.24U L=0.12U M=1 
X2 net28 A VSS VSS LPNFET W=1.38U L=0.12U M=1 
X3 net28 nmen VSS VSS LPNFET W=0.46U L=0.12U M=1 
X4 Y net28 VSS VSS LPNFET W=3.5U L=0.12U M=1 
X5 nmin OE net28 VSS LPNFET W=0.74U L=0.12U M=1 
X6 nmin A VDD VDD LPPFET W=2.06U L=0.12U M=1 
X7 nmin OE VDD VDD LPPFET W=0.62U L=0.12U M=1 
X8 net28 nmen nmin VDD LPPFET W=1.02U L=0.12U M=1 
X9 Y nmin VDD VDD LPPFET W=4.98U L=0.12U M=1 
.ENDS TBUFX8TS 

**** 
*.SUBCKT TBUFXLTS Y A OE 
.SUBCKT TBUFXLTS Y A OE VSS VDD
X0 VDD OE nmen VDD LPPFET W=0.28U L=0.12U M=1 
X1 nmen OE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 net28 A VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 net28 nmen VSS VSS LPNFET W=0.18U L=0.12U M=1 
X4 Y net28 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X5 nmin OE net28 VSS LPNFET W=0.2U L=0.12U M=1 
X6 nmin A VDD VDD LPPFET W=0.28U L=0.12U M=1 
X7 nmin OE VDD VDD LPPFET W=0.28U L=0.12U M=1 
X8 net28 nmen nmin VDD LPPFET W=0.28U L=0.12U M=1 
X9 Y nmin VDD VDD LPPFET W=0.42U L=0.12U M=1 
.ENDS TBUFXLTS 

**** 
*.SUBCKT TIEHITS Y 
.SUBCKT TIEHITS Y VSS VDD
X0 net4 net4 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X1 Y net4 VDD VDD LPPFET W=0.64U L=0.12U M=1 
.ENDS TIEHITS 

**** 
*.SUBCKT TIELOTS Y 
.SUBCKT TIELOTS Y VSS VDD
X0 Y net7 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X1 net7 net7 VDD VDD LPPFET W=0.28U L=0.12U M=1 
.ENDS TIELOTS 

**** 
*.SUBCKT TLATNCAX12TS ECK CK E 
.SUBCKT TLATNCAX12TS ECK CK E VSS VDD
X0 net23 c VSS VSS LPNFET W=0.44U L=0.12U M=1 
X1 net23 nmin VSS VSS LPNFET W=0.44U L=0.12U M=1 
X10 hnet27 c nmin VDD LPPFET W=0.28U L=0.12U M=1 
X11 VDD m hnet27 VDD LPPFET W=0.28U L=0.12U M=1 
X12 VDD net35 ECK VDD LPPFET W=14.3U L=0.12U M=1 
X13 ECK net35 VSS VSS LPNFET W=5.52U L=0.12U M=1 
X14 VDD net23 net35 VDD LPPFET W=4.76U L=0.12U M=1 
X15 net35 net23 VSS VSS LPNFET W=1.8U L=0.12U M=1 
X16 VDD c cn VDD LPPFET W=0.28U L=0.12U M=1 
X17 cn c VSS VSS LPNFET W=0.2U L=0.12U M=1 
X18 VDD CK c VDD LPPFET W=0.84U L=0.12U M=1 
X19 c CK VSS VSS LPNFET W=0.6U L=0.12U M=1 
X2 VDD c hnet13 VDD LPPFET W=1.3U L=0.12U M=1 
X20 VDD nmin m VDD LPPFET W=0.28U L=0.12U M=1 
X21 m nmin VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 hnet13 nmin net23 VDD LPPFET W=1.3U L=0.12U M=1 
X4 hnet19 E VSS VSS LPNFET W=0.82U L=0.12U M=1 
X5 nmin c hnet19 VSS LPNFET W=0.82U L=0.12U M=1 
X6 hnet21 cn nmin VDD LPPFET W=1.14U L=0.12U M=1 
X7 VDD E hnet21 VDD LPPFET W=1.14U L=0.12U M=1 
X8 hnet25 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X9 nmin cn hnet25 VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS TLATNCAX12TS 

**** 
*.SUBCKT TLATNCAX16TS ECK CK E 
.SUBCKT TLATNCAX16TS ECK CK E VSS VDD
X0 net23 c VSS VSS LPNFET W=0.58U L=0.12U M=1 
X1 net23 nmin VSS VSS LPNFET W=0.58U L=0.12U M=1 
X10 hnet26 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X11 nmin cn hnet26 VSS LPNFET W=0.2U L=0.12U M=1 
X12 hnet28 c nmin VDD LPPFET W=0.28U L=0.12U M=1 
X13 VDD m hnet28 VDD LPPFET W=0.28U L=0.12U M=1 
X14 VDD net35 ECK VDD LPPFET W=18.9U L=0.12U M=1 
X15 ECK net35 VSS VSS LPNFET W=7.36U L=0.12U M=1 
X16 VDD net23 net35 VDD LPPFET W=6.3U L=0.12U M=1 
X17 net35 net23 VSS VSS LPNFET W=2.34U L=0.12U M=1 
X18 VDD c cn VDD LPPFET W=0.3U L=0.12U M=1 
X19 cn c VSS VSS LPNFET W=0.22U L=0.12U M=1 
X2 VDD c hnet14 VDD LPPFET W=0.98U L=0.12U M=1 
X20 VDD CK c VDD LPPFET W=1.02U L=0.12U M=1 
X21 c CK VSS VSS LPNFET W=0.74U L=0.12U M=1 
X22 VDD nmin m VDD LPPFET W=0.28U L=0.12U M=1 
X23 m nmin VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 hnet14 nmin net23 VDD LPPFET W=0.98U L=0.12U M=1 
X4 VDD c hnet12 VDD LPPFET W=0.98U L=0.12U M=1 
X5 hnet12 nmin net23 VDD LPPFET W=0.98U L=0.12U M=1 
X6 hnet20 E VSS VSS LPNFET W=0.84U L=0.12U M=1 
X7 nmin c hnet20 VSS LPNFET W=0.84U L=0.12U M=1 
X8 hnet22 cn nmin VDD LPPFET W=1.26U L=0.12U M=1 
X9 VDD E hnet22 VDD LPPFET W=1.26U L=0.12U M=1 
.ENDS TLATNCAX16TS 

**** 
*.SUBCKT TLATNCAX20TS ECK CK E 
.SUBCKT TLATNCAX20TS ECK CK E VSS VDD
X0 net23 c VSS VSS LPNFET W=0.74U L=0.12U M=1 
X1 net23 nmin VSS VSS LPNFET W=0.74U L=0.12U M=1 
X10 hnet26 cn nmin VDD LPPFET W=0.88U L=0.12U M=1 
X11 hnet24 cn nmin VDD LPPFET W=0.88U L=0.12U M=1 
X12 VDD E hnet26 VDD LPPFET W=0.88U L=0.12U M=1 
X13 VDD E hnet24 VDD LPPFET W=0.88U L=0.12U M=1 
X14 hnet28 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X15 nmin cn hnet28 VSS LPNFET W=0.2U L=0.12U M=1 
X16 hnet30 c nmin VDD LPPFET W=0.28U L=0.12U M=1 
X17 VDD m hnet30 VDD LPPFET W=0.28U L=0.12U M=1 
X18 VDD net36 ECK VDD LPPFET W=21.6U L=0.12U M=1 
X19 ECK net36 VSS VSS LPNFET W=8.28U L=0.12U M=1 
X2 VDD c hnet14 VDD LPPFET W=1.3U L=0.12U M=1 
X20 VDD net23 net36 VDD LPPFET W=7.8U L=0.12U M=1 
X21 net36 net23 VSS VSS LPNFET W=2.94U L=0.12U M=1 
X22 VDD c cn VDD LPPFET W=0.42U L=0.12U M=1 
X23 cn c VSS VSS LPNFET W=0.3U L=0.12U M=1 
X24 VDD CK c VDD LPPFET W=1.3U L=0.12U M=1 
X25 c CK VSS VSS LPNFET W=0.92U L=0.12U M=1 
X26 VDD nmin m VDD LPPFET W=0.28U L=0.12U M=1 
X27 m nmin VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 hnet14 nmin net23 VDD LPPFET W=1.3U L=0.12U M=1 
X4 VDD c hnet12 VDD LPPFET W=1.3U L=0.12U M=1 
X5 hnet12 nmin net23 VDD LPPFET W=1.3U L=0.12U M=1 
X6 hnet20 E VSS VSS LPNFET W=0.6U L=0.12U M=1 
X7 hnet21 E VSS VSS LPNFET W=0.6U L=0.12U M=1 
X8 nmin c hnet20 VSS LPNFET W=0.6U L=0.12U M=1 
X9 nmin c hnet21 VSS LPNFET W=0.6U L=0.12U M=1 
.ENDS TLATNCAX20TS 

**** 
*.SUBCKT TLATNCAX2TS ECK CK E 
.SUBCKT TLATNCAX2TS ECK CK E VSS VDD
X0 ECK c VSS VSS LPNFET W=0.38U L=0.12U M=1 
X1 ECK nmin VSS VSS LPNFET W=0.38U L=0.12U M=1 
X10 hnet25 c nmin VDD LPPFET W=0.28U L=0.12U M=1 
X11 VDD m hnet25 VDD LPPFET W=0.28U L=0.12U M=1 
X12 VDD c cn VDD LPPFET W=0.28U L=0.12U M=1 
X13 cn c VSS VSS LPNFET W=0.2U L=0.12U M=1 
X14 VDD CK c VDD LPPFET W=0.72U L=0.12U M=1 
X15 c CK VSS VSS LPNFET W=0.52U L=0.12U M=1 
X16 VDD nmin m VDD LPPFET W=0.28U L=0.12U M=1 
X17 m nmin VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 VDD c hnet11 VDD LPPFET W=1.3U L=0.12U M=1 
X3 hnet11 nmin ECK VDD LPPFET W=1.3U L=0.12U M=1 
X4 hnet17 E VSS VSS LPNFET W=0.72U L=0.12U M=1 
X5 nmin c hnet17 VSS LPNFET W=0.72U L=0.12U M=1 
X6 hnet19 cn nmin VDD LPPFET W=1U L=0.12U M=1 
X7 VDD E hnet19 VDD LPPFET W=1U L=0.12U M=1 
X8 hnet23 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X9 nmin cn hnet23 VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS TLATNCAX2TS 

**** 
*.SUBCKT TLATNCAX3TS ECK CK E 
.SUBCKT TLATNCAX3TS ECK CK E VSS VDD
X0 ECK c VSS VSS LPNFET W=0.56U L=0.12U M=1 
X1 ECK nmin VSS VSS LPNFET W=0.56U L=0.12U M=1 
X10 hnet24 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X11 nmin cn hnet24 VSS LPNFET W=0.2U L=0.12U M=1 
X12 hnet26 c nmin VDD LPPFET W=0.28U L=0.12U M=1 
X13 VDD m hnet26 VDD LPPFET W=0.28U L=0.12U M=1 
X14 VDD c cn VDD LPPFET W=0.3U L=0.12U M=1 
X15 cn c VSS VSS LPNFET W=0.22U L=0.12U M=1 
X16 VDD CK c VDD LPPFET W=1U L=0.12U M=1 
X17 c CK VSS VSS LPNFET W=0.72U L=0.12U M=1 
X18 VDD nmin m VDD LPPFET W=0.28U L=0.12U M=1 
X19 m nmin VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 VDD c hnet12 VDD LPPFET W=0.96U L=0.12U M=1 
X3 hnet12 nmin ECK VDD LPPFET W=0.96U L=0.12U M=1 
X4 VDD c hnet10 VDD LPPFET W=0.96U L=0.12U M=1 
X5 hnet10 nmin ECK VDD LPPFET W=0.96U L=0.12U M=1 
X6 hnet18 E VSS VSS LPNFET W=0.82U L=0.12U M=1 
X7 nmin c hnet18 VSS LPNFET W=0.82U L=0.12U M=1 
X8 hnet20 cn nmin VDD LPPFET W=1.26U L=0.12U M=1 
X9 VDD E hnet20 VDD LPPFET W=1.26U L=0.12U M=1 
.ENDS TLATNCAX3TS 

**** 
*.SUBCKT TLATNCAX4TS ECK CK E 
.SUBCKT TLATNCAX4TS ECK CK E VSS VDD
X0 ECK c VSS VSS LPNFET W=0.74U L=0.12U M=1 
X1 ECK nmin VSS VSS LPNFET W=0.74U L=0.12U M=1 
X10 hnet24 cn nmin VDD LPPFET W=0.88U L=0.12U M=1 
X11 hnet22 cn nmin VDD LPPFET W=0.88U L=0.12U M=1 
X12 VDD E hnet24 VDD LPPFET W=0.88U L=0.12U M=1 
X13 VDD E hnet22 VDD LPPFET W=0.88U L=0.12U M=1 
X14 hnet26 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X15 nmin cn hnet26 VSS LPNFET W=0.2U L=0.12U M=1 
X16 hnet28 c nmin VDD LPPFET W=0.28U L=0.12U M=1 
X17 VDD m hnet28 VDD LPPFET W=0.28U L=0.12U M=1 
X18 VDD c cn VDD LPPFET W=0.42U L=0.12U M=1 
X19 cn c VSS VSS LPNFET W=0.3U L=0.12U M=1 
X2 VDD c hnet12 VDD LPPFET W=1.28U L=0.12U M=1 
X20 VDD CK c VDD LPPFET W=1.3U L=0.12U M=1 
X21 c CK VSS VSS LPNFET W=0.92U L=0.12U M=1 
X22 VDD nmin m VDD LPPFET W=0.28U L=0.12U M=1 
X23 m nmin VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 hnet12 nmin ECK VDD LPPFET W=1.28U L=0.12U M=1 
X4 VDD c hnet10 VDD LPPFET W=1.28U L=0.12U M=1 
X5 hnet10 nmin ECK VDD LPPFET W=1.28U L=0.12U M=1 
X6 hnet18 E VSS VSS LPNFET W=0.6U L=0.12U M=1 
X7 hnet19 E VSS VSS LPNFET W=0.6U L=0.12U M=1 
X8 nmin c hnet18 VSS LPNFET W=0.6U L=0.12U M=1 
X9 nmin c hnet19 VSS LPNFET W=0.6U L=0.12U M=1 
.ENDS TLATNCAX4TS 

**** 
*.SUBCKT TLATNCAX6TS ECK CK E 
.SUBCKT TLATNCAX6TS ECK CK E VSS VDD
X0 ECK c VSS VSS LPNFET W=1.12U L=0.12U M=1 
X1 ECK nmin VSS VSS LPNFET W=1.12U L=0.12U M=1 
X10 nmin c hnet19 VSS LPNFET W=0.88U L=0.12U M=1 
X11 nmin c hnet20 VSS LPNFET W=0.88U L=0.12U M=1 
X12 hnet25 cn nmin VDD LPPFET W=1.22U L=0.12U M=1 
X13 hnet23 cn nmin VDD LPPFET W=1.22U L=0.12U M=1 
X14 VDD E hnet25 VDD LPPFET W=1.22U L=0.12U M=1 
X15 VDD E hnet23 VDD LPPFET W=1.22U L=0.12U M=1 
X16 hnet27 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X17 nmin cn hnet27 VSS LPNFET W=0.2U L=0.12U M=1 
X18 hnet29 c nmin VDD LPPFET W=0.28U L=0.12U M=1 
X19 VDD m hnet29 VDD LPPFET W=0.28U L=0.12U M=1 
X2 VDD c hnet12 VDD LPPFET W=1.28U L=0.12U M=1 
X20 VDD c cn VDD LPPFET W=0.56U L=0.12U M=1 
X21 cn c VSS VSS LPNFET W=0.4U L=0.12U M=1 
X22 VDD CK c VDD LPPFET W=1.92U L=0.12U M=1 
X23 c CK VSS VSS LPNFET W=1.32U L=0.12U M=1 
X24 VDD nmin m VDD LPPFET W=0.28U L=0.12U M=1 
X25 m nmin VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 hnet12 nmin ECK VDD LPPFET W=1.28U L=0.12U M=1 
X4 VDD c hnet10 VDD LPPFET W=1.28U L=0.12U M=1 
X5 hnet10 nmin ECK VDD LPPFET W=1.28U L=0.12U M=1 
X6 VDD c hnet14 VDD LPPFET W=1.28U L=0.12U M=1 
X7 hnet14 nmin ECK VDD LPPFET W=1.28U L=0.12U M=1 
X8 hnet19 E VSS VSS LPNFET W=0.88U L=0.12U M=1 
X9 hnet20 E VSS VSS LPNFET W=0.88U L=0.12U M=1 
.ENDS TLATNCAX6TS 

**** 
*.SUBCKT TLATNCAX8TS ECK CK E 
.SUBCKT TLATNCAX8TS ECK CK E VSS VDD
X0 ECK c VSS VSS LPNFET W=1.86U L=0.12U M=1 
X1 ECK nmin VSS VSS LPNFET W=1.86U L=0.12U M=1 
X10 VDD c hnet13 VDD LPPFET W=1.3U L=0.12U M=1 
X11 hnet13 nmin ECK VDD LPPFET W=1.3U L=0.12U M=1 
X12 VDD c hnet10 VDD LPPFET W=1.3U L=0.12U M=1 
X13 hnet10 nmin ECK VDD LPPFET W=1.3U L=0.12U M=1 
X14 VDD c hnet20 VDD LPPFET W=1.3U L=0.12U M=1 
X15 hnet20 nmin ECK VDD LPPFET W=1.3U L=0.12U M=1 
X16 hnet23 E VSS VSS LPNFET W=0.84U L=0.12U M=1 
X17 hnet25 E VSS VSS LPNFET W=0.84U L=0.12U M=1 
X18 hnet32 E VSS VSS LPNFET W=0.84U L=0.12U M=1 
X19 hnet24 E VSS VSS LPNFET W=0.84U L=0.12U M=1 
X2 VDD c hnet17 VDD LPPFET W=1.3U L=0.12U M=1 
X20 nmin c hnet23 VSS LPNFET W=0.84U L=0.12U M=1 
X21 nmin c hnet25 VSS LPNFET W=0.84U L=0.12U M=1 
X22 nmin c hnet32 VSS LPNFET W=0.84U L=0.12U M=1 
X23 nmin c hnet24 VSS LPNFET W=0.84U L=0.12U M=1 
X24 hnet30 cn nmin VDD LPPFET W=1.26U L=0.12U M=1 
X25 hnet33 cn nmin VDD LPPFET W=1.26U L=0.12U M=1 
X26 hnet26 cn nmin VDD LPPFET W=1.26U L=0.12U M=1 
X27 hnet31 cn nmin VDD LPPFET W=1.26U L=0.12U M=1 
X28 VDD E hnet30 VDD LPPFET W=1.26U L=0.12U M=1 
X29 VDD E hnet33 VDD LPPFET W=1.26U L=0.12U M=1 
X3 hnet17 nmin ECK VDD LPPFET W=1.3U L=0.12U M=1 
X30 VDD E hnet26 VDD LPPFET W=1.26U L=0.12U M=1 
X31 VDD E hnet31 VDD LPPFET W=1.26U L=0.12U M=1 
X32 hnet35 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X33 nmin cn hnet35 VSS LPNFET W=0.2U L=0.12U M=1 
X34 hnet37 c nmin VDD LPPFET W=0.28U L=0.12U M=1 
X35 VDD m hnet37 VDD LPPFET W=0.28U L=0.12U M=1 
X36 VDD c cn VDD LPPFET W=1.08U L=0.12U M=1 
X37 cn c VSS VSS LPNFET W=0.78U L=0.12U M=1 
X38 VDD CK c VDD LPPFET W=3.9U L=0.12U M=1 
X39 c CK VSS VSS LPNFET W=2.76U L=0.12U M=1 
X4 VDD c hnet11 VDD LPPFET W=1.3U L=0.12U M=1 
X40 VDD nmin m VDD LPPFET W=0.28U L=0.12U M=1 
X41 m nmin VSS VSS LPNFET W=0.2U L=0.12U M=1 
X5 hnet11 nmin ECK VDD LPPFET W=1.3U L=0.12U M=1 
X6 VDD c hnet16 VDD LPPFET W=1.3U L=0.12U M=1 
X7 hnet16 nmin ECK VDD LPPFET W=1.3U L=0.12U M=1 
X8 VDD c hnet15 VDD LPPFET W=1.3U L=0.12U M=1 
X9 hnet15 nmin ECK VDD LPPFET W=1.3U L=0.12U M=1 
.ENDS TLATNCAX8TS 

**** 
*.SUBCKT TLATNSRX1TS Q QN D GN RN SN 
.SUBCKT TLATNSRX1TS Q QN D GN RN SN VSS VDD
X0 VDD D hnet20 VDD LPPFET W=0.54U L=0.12U M=1 
X1 hnet20 nms hnet25 VDD LPPFET W=0.54U L=0.12U M=1 
X10 VDD pm Q VDD LPPFET W=0.58U L=0.12U M=1 
X11 Q pm VSS VSS LPNFET W=0.42U L=0.12U M=1 
X12 VDD SN nms VDD LPPFET W=0.42U L=0.12U M=1 
X13 nms SN VSS VSS LPNFET W=0.3U L=0.12U M=1 
X14 VDD c cn VDD LPPFET W=0.28U L=0.12U M=1 
X15 cn c VSS VSS LPNFET W=0.2U L=0.12U M=1 
X16 VDD GN c VDD LPPFET W=0.38U L=0.12U M=1 
X17 c GN VSS VSS LPNFET W=0.26U L=0.12U M=1 
X18 VDD pm m VDD LPPFET W=0.3U L=0.12U M=1 
X19 m pm VSS VSS LPNFET W=0.22U L=0.12U M=1 
X2 hnet25 cn pm VDD LPPFET W=0.54U L=0.12U M=1 
X20 net66 nms net72 VDD LPPFET W=0.36U L=0.12U M=1 
X21 pm c net66 VDD LPPFET W=0.36U L=0.12U M=1 
X22 net72 m VDD VDD LPPFET W=0.36U L=0.12U M=1 
X23 net75 RN net78 VSS LPNFET W=0.32U L=0.12U M=1 
X24 net78 m VSS VSS LPNFET W=0.32U L=0.12U M=1 
X25 pm cn net75 VSS LPNFET W=0.32U L=0.12U M=1 
X26 pm nms VSS VSS LPNFET W=0.28U L=0.12U M=1 
X3 hnet31 D VSS VSS LPNFET W=0.42U L=0.12U M=1 
X4 hnet26 RN hnet31 VSS LPNFET W=0.42U L=0.12U M=1 
X5 pm c hnet26 VSS LPNFET W=0.42U L=0.12U M=1 
X6 VDD RN hnet35 VDD LPPFET W=0.48U L=0.12U M=1 
X7 hnet35 nms pm VDD LPPFET W=0.48U L=0.12U M=1 
X8 VDD m QN VDD LPPFET W=0.54U L=0.12U M=1 
X9 QN m VSS VSS LPNFET W=0.46U L=0.12U M=1 
.ENDS TLATNSRX1TS 

**** 
*.SUBCKT TLATNSRX2TS Q QN D GN RN SN 
.SUBCKT TLATNSRX2TS Q QN D GN RN SN VSS VDD
X0 VDD D hnet20 VDD LPPFET W=1.12U L=0.12U M=1 
X1 hnet20 nms hnet25 VDD LPPFET W=1.12U L=0.12U M=1 
X10 VDD pm Q VDD LPPFET W=1.28U L=0.12U M=1 
X11 Q pm VSS VSS LPNFET W=0.9U L=0.12U M=1 
X12 VDD SN nms VDD LPPFET W=0.66U L=0.12U M=1 
X13 nms SN VSS VSS LPNFET W=0.48U L=0.12U M=1 
X14 VDD c cn VDD LPPFET W=0.28U L=0.12U M=1 
X15 cn c VSS VSS LPNFET W=0.22U L=0.12U M=1 
X16 VDD GN c VDD LPPFET W=0.42U L=0.12U M=1 
X17 c GN VSS VSS LPNFET W=0.3U L=0.12U M=1 
X18 VDD pm m VDD LPPFET W=0.48U L=0.12U M=1 
X19 m pm VSS VSS LPNFET W=0.34U L=0.12U M=1 
X2 hnet25 cn pm VDD LPPFET W=1.12U L=0.12U M=1 
X20 net66 nms net72 VDD LPPFET W=0.36U L=0.12U M=1 
X21 pm c net66 VDD LPPFET W=0.36U L=0.12U M=1 
X22 net72 m VDD VDD LPPFET W=0.36U L=0.12U M=1 
X23 net75 RN net78 VSS LPNFET W=0.32U L=0.12U M=1 
X24 net78 m VSS VSS LPNFET W=0.32U L=0.12U M=1 
X25 pm cn net75 VSS LPNFET W=0.32U L=0.12U M=1 
X26 pm nms VSS VSS LPNFET W=0.5U L=0.12U M=1 
X3 hnet31 D VSS VSS LPNFET W=0.74U L=0.12U M=1 
X4 hnet26 RN hnet31 VSS LPNFET W=0.74U L=0.12U M=1 
X5 pm c hnet26 VSS LPNFET W=0.74U L=0.12U M=1 
X6 VDD RN hnet35 VDD LPPFET W=0.92U L=0.12U M=1 
X7 hnet35 nms pm VDD LPPFET W=0.92U L=0.12U M=1 
X8 VDD m QN VDD LPPFET W=1.28U L=0.12U M=1 
X9 QN m VSS VSS LPNFET W=0.9U L=0.12U M=1 
.ENDS TLATNSRX2TS 

**** 
*.SUBCKT TLATNSRX4TS Q QN D GN RN SN 
.SUBCKT TLATNSRX4TS Q QN D GN RN SN VSS VDD
X0 hnet27 D VSS VSS LPNFET W=0.48U L=0.12U M=1 
X1 hnet20 RN hnet27 VSS LPNFET W=0.48U L=0.12U M=1 
X10 hnet31 nms hnet30 VDD LPPFET W=0.98U L=0.12U M=1 
X11 hnet30 cn pm VDD LPPFET W=0.98U L=0.12U M=1 
X12 VDD D hnet33 VDD LPPFET W=0.98U L=0.12U M=1 
X13 hnet33 nms hnet34 VDD LPPFET W=0.98U L=0.12U M=1 
X14 hnet34 cn pm VDD LPPFET W=0.98U L=0.12U M=1 
X15 VDD RN hnet42 VDD LPPFET W=0.92U L=0.12U M=1 
X16 hnet42 nms pm VDD LPPFET W=0.92U L=0.12U M=1 
X17 VDD RN hnet39 VDD LPPFET W=0.92U L=0.12U M=1 
X18 hnet39 nms pm VDD LPPFET W=0.92U L=0.12U M=1 
X19 VDD m QN VDD LPPFET W=2.56U L=0.12U M=1 
X2 pm c hnet20 VSS LPNFET W=0.48U L=0.12U M=1 
X20 QN m VSS VSS LPNFET W=1.84U L=0.12U M=1 
X21 VDD pm Q VDD LPPFET W=2.56U L=0.12U M=1 
X22 Q pm VSS VSS LPNFET W=1.84U L=0.12U M=1 
X23 VDD SN nms VDD LPPFET W=1.22U L=0.12U M=1 
X24 nms SN VSS VSS LPNFET W=0.88U L=0.12U M=1 
X25 VDD c cn VDD LPPFET W=0.5U L=0.12U M=1 
X26 cn c VSS VSS LPNFET W=0.36U L=0.12U M=1 
X27 VDD GN c VDD LPPFET W=0.7U L=0.12U M=1 
X28 c GN VSS VSS LPNFET W=0.5U L=0.12U M=1 
X29 VDD pm m VDD LPPFET W=0.84U L=0.12U M=1 
X3 hnet29 D VSS VSS LPNFET W=0.48U L=0.12U M=1 
X30 m pm VSS VSS LPNFET W=0.6U L=0.12U M=1 
X31 net66 nms net72 VDD LPPFET W=0.32U L=0.12U M=1 
X32 pm c net66 VDD LPPFET W=0.32U L=0.12U M=1 
X33 net72 m VDD VDD LPPFET W=0.32U L=0.12U M=1 
X34 net75 RN net78 VSS LPNFET W=0.32U L=0.12U M=1 
X35 net78 m VSS VSS LPNFET W=0.32U L=0.12U M=1 
X36 pm cn net75 VSS LPNFET W=0.32U L=0.12U M=1 
X37 pm nms VSS VSS LPNFET W=0.92U L=0.12U M=1 
X4 hnet28 RN hnet29 VSS LPNFET W=0.48U L=0.12U M=1 
X5 pm c hnet28 VSS LPNFET W=0.48U L=0.12U M=1 
X6 hnet23 D VSS VSS LPNFET W=0.48U L=0.12U M=1 
X7 hnet21 RN hnet23 VSS LPNFET W=0.48U L=0.12U M=1 
X8 pm c hnet21 VSS LPNFET W=0.48U L=0.12U M=1 
X9 VDD D hnet31 VDD LPPFET W=0.98U L=0.12U M=1 
.ENDS TLATNSRX4TS 

**** 
*.SUBCKT TLATNSRXLTS Q QN D GN RN SN 
.SUBCKT TLATNSRXLTS Q QN D GN RN SN VSS VDD
X0 VDD D hnet20 VDD LPPFET W=0.36U L=0.12U M=1 
X1 hnet20 nms hnet25 VDD LPPFET W=0.36U L=0.12U M=1 
X10 VDD pm Q VDD LPPFET W=0.42U L=0.12U M=1 
X11 Q pm VSS VSS LPNFET W=0.24U L=0.12U M=1 
X12 VDD SN nms VDD LPPFET W=0.28U L=0.12U M=1 
X13 nms SN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X14 VDD c cn VDD LPPFET W=0.28U L=0.12U M=1 
X15 cn c VSS VSS LPNFET W=0.2U L=0.12U M=1 
X16 VDD GN c VDD LPPFET W=0.28U L=0.12U M=1 
X17 c GN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X18 VDD pm m VDD LPPFET W=0.28U L=0.12U M=1 
X19 m pm VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 hnet25 cn pm VDD LPPFET W=0.36U L=0.12U M=1 
X20 net66 nms net72 VDD LPPFET W=0.36U L=0.12U M=1 
X21 pm c net66 VDD LPPFET W=0.36U L=0.12U M=1 
X22 net72 m VDD VDD LPPFET W=0.36U L=0.12U M=1 
X23 net75 RN net78 VSS LPNFET W=0.32U L=0.12U M=1 
X24 net78 m VSS VSS LPNFET W=0.32U L=0.12U M=1 
X25 pm cn net75 VSS LPNFET W=0.32U L=0.12U M=1 
X26 pm nms VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 hnet31 D VSS VSS LPNFET W=0.32U L=0.12U M=1 
X4 hnet26 RN hnet31 VSS LPNFET W=0.32U L=0.12U M=1 
X5 pm c hnet26 VSS LPNFET W=0.32U L=0.12U M=1 
X6 VDD RN hnet35 VDD LPPFET W=0.3U L=0.12U M=1 
X7 hnet35 nms pm VDD LPPFET W=0.3U L=0.12U M=1 
X8 VDD m QN VDD LPPFET W=0.42U L=0.12U M=1 
X9 QN m VSS VSS LPNFET W=0.24U L=0.12U M=1 
.ENDS TLATNSRXLTS 

**** 
*.SUBCKT TLATNTSCAX12TS ECK CK E SE 
.SUBCKT TLATNTSCAX12TS ECK CK E SE VSS VDD
X0 net27 SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X1 net27 E VSS VSS LPNFET W=0.2U L=0.12U M=1 
X10 hnet30 cn net34 VDD LPPFET W=1.14U L=0.12U M=1 
X11 VDD net45 hnet30 VDD LPPFET W=1.14U L=0.12U M=1 
X12 hnet34 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X13 net34 cn hnet34 VSS LPNFET W=0.2U L=0.12U M=1 
X14 hnet36 c net34 VDD LPPFET W=0.28U L=0.12U M=1 
X15 VDD m hnet36 VDD LPPFET W=0.28U L=0.12U M=1 
X16 VDD net43 ECK VDD LPPFET W=14.9U L=0.12U M=1 
X17 ECK net43 VSS VSS LPNFET W=5.48U L=0.12U M=1 
X18 VDD net30 net43 VDD LPPFET W=4.28U L=0.12U M=1 
X19 net43 net30 VSS VSS LPNFET W=1.58U L=0.12U M=1 
X2 VDD SE hnet16 VDD LPPFET W=0.36U L=0.12U M=1 
X20 VDD net27 net45 VDD LPPFET W=0.44U L=0.12U M=1 
X21 net45 net27 VSS VSS LPNFET W=0.32U L=0.12U M=1 
X22 VDD c cn VDD LPPFET W=0.28U L=0.12U M=1 
X23 cn c VSS VSS LPNFET W=0.2U L=0.12U M=1 
X24 VDD CK c VDD LPPFET W=0.84U L=0.12U M=1 
X25 c CK VSS VSS LPNFET W=0.6U L=0.12U M=1 
X26 VDD net34 m VDD LPPFET W=0.28U L=0.12U M=1 
X27 m net34 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 hnet16 E net27 VDD LPPFET W=0.36U L=0.12U M=1 
X4 net30 c VSS VSS LPNFET W=0.44U L=0.12U M=1 
X5 net30 net34 VSS VSS LPNFET W=0.44U L=0.12U M=1 
X6 VDD c hnet22 VDD LPPFET W=1.42U L=0.12U M=1 
X7 hnet22 net34 net30 VDD LPPFET W=1.42U L=0.12U M=1 
X8 hnet28 net45 VSS VSS LPNFET W=0.82U L=0.12U M=1 
X9 net34 c hnet28 VSS LPNFET W=0.82U L=0.12U M=1 
.ENDS TLATNTSCAX12TS 

**** 
*.SUBCKT TLATNTSCAX16TS ECK CK E SE 
.SUBCKT TLATNTSCAX16TS ECK CK E SE VSS VDD
X0 net27 SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X1 net27 E VSS VSS LPNFET W=0.2U L=0.12U M=1 
X10 hnet27 net45 VSS VSS LPNFET W=0.84U L=0.12U M=1 
X11 net34 c hnet27 VSS LPNFET W=0.84U L=0.12U M=1 
X12 hnet29 cn net34 VDD LPPFET W=1.28U L=0.12U M=1 
X13 VDD net45 hnet29 VDD LPPFET W=1.28U L=0.12U M=1 
X14 hnet33 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X15 net34 cn hnet33 VSS LPNFET W=0.2U L=0.12U M=1 
X16 hnet35 c net34 VDD LPPFET W=0.28U L=0.12U M=1 
X17 VDD m hnet35 VDD LPPFET W=0.28U L=0.12U M=1 
X18 VDD net43 ECK VDD LPPFET W=19.86U L=0.12U M=1 
X19 ECK net43 VSS VSS LPNFET W=7.36U L=0.12U M=1 
X2 VDD SE hnet16 VDD LPPFET W=0.36U L=0.12U M=1 
X20 VDD net30 net43 VDD LPPFET W=5.68U L=0.12U M=1 
X21 net43 net30 VSS VSS LPNFET W=2.32U L=0.12U M=1 
X22 VDD net27 net45 VDD LPPFET W=0.5U L=0.12U M=1 
X23 net45 net27 VSS VSS LPNFET W=0.36U L=0.12U M=1 
X24 VDD c cn VDD LPPFET W=0.3U L=0.12U M=1 
X25 cn c VSS VSS LPNFET W=0.22U L=0.12U M=1 
X26 VDD CK c VDD LPPFET W=1.02U L=0.12U M=1 
X27 c CK VSS VSS LPNFET W=0.74U L=0.12U M=1 
X28 VDD net34 m VDD LPPFET W=0.28U L=0.12U M=1 
X29 m net34 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 hnet16 E net27 VDD LPPFET W=0.36U L=0.12U M=1 
X4 net30 c VSS VSS LPNFET W=0.58U L=0.12U M=1 
X5 net30 net34 VSS VSS LPNFET W=0.58U L=0.12U M=1 
X6 VDD c hnet23 VDD LPPFET W=1U L=0.12U M=1 
X7 hnet23 net34 net30 VDD LPPFET W=1U L=0.12U M=1 
X8 VDD c hnet21 VDD LPPFET W=1U L=0.12U M=1 
X9 hnet21 net34 net30 VDD LPPFET W=1U L=0.12U M=1 
.ENDS TLATNTSCAX16TS 

**** 
*.SUBCKT TLATNTSCAX20TS ECK CK E SE 
.SUBCKT TLATNTSCAX20TS ECK CK E SE VSS VDD
X0 net27 SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X1 net27 E VSS VSS LPNFET W=0.2U L=0.12U M=1 
X10 hnet27 net45 VSS VSS LPNFET W=0.64U L=0.12U M=1 
X11 hnet28 net45 VSS VSS LPNFET W=0.64U L=0.12U M=1 
X12 net34 c hnet27 VSS LPNFET W=0.64U L=0.12U M=1 
X13 net34 c hnet28 VSS LPNFET W=0.64U L=0.12U M=1 
X14 hnet33 cn net34 VDD LPPFET W=0.86U L=0.12U M=1 
X15 hnet31 cn net34 VDD LPPFET W=0.86U L=0.12U M=1 
X16 VDD net45 hnet33 VDD LPPFET W=0.86U L=0.12U M=1 
X17 VDD net45 hnet31 VDD LPPFET W=0.86U L=0.12U M=1 
X18 hnet35 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X19 net34 cn hnet35 VSS LPNFET W=0.2U L=0.12U M=1 
X2 VDD SE hnet16 VDD LPPFET W=0.36U L=0.12U M=1 
X20 hnet37 c net34 VDD LPPFET W=0.28U L=0.12U M=1 
X21 VDD m hnet37 VDD LPPFET W=0.28U L=0.12U M=1 
X22 VDD net42 ECK VDD LPPFET W=23.36U L=0.12U M=1 
X23 ECK net42 VSS VSS LPNFET W=9.2U L=0.12U M=1 
X24 VDD net30 net42 VDD LPPFET W=8.04U L=0.12U M=1 
X25 net42 net30 VSS VSS LPNFET W=2.94U L=0.12U M=1 
X26 VDD net27 net45 VDD LPPFET W=0.7U L=0.12U M=1 
X27 net45 net27 VSS VSS LPNFET W=0.5U L=0.12U M=1 
X28 VDD c cn VDD LPPFET W=0.42U L=0.12U M=1 
X29 cn c VSS VSS LPNFET W=0.3U L=0.12U M=1 
X3 hnet16 E net27 VDD LPPFET W=0.36U L=0.12U M=1 
X30 VDD CK c VDD LPPFET W=1.36U L=0.12U M=1 
X31 c CK VSS VSS LPNFET W=0.92U L=0.12U M=1 
X32 VDD net34 m VDD LPPFET W=0.28U L=0.12U M=1 
X33 m net34 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X4 net30 c VSS VSS LPNFET W=0.74U L=0.12U M=1 
X5 net30 net34 VSS VSS LPNFET W=0.74U L=0.12U M=1 
X6 VDD c hnet23 VDD LPPFET W=1.28U L=0.12U M=1 
X7 hnet23 net34 net30 VDD LPPFET W=1.28U L=0.12U M=1 
X8 VDD c hnet21 VDD LPPFET W=1.28U L=0.12U M=1 
X9 hnet21 net34 net30 VDD LPPFET W=1.28U L=0.12U M=1 
.ENDS TLATNTSCAX20TS 

**** 
*.SUBCKT TLATNTSCAX2TS ECK CK E SE 
.SUBCKT TLATNTSCAX2TS ECK CK E SE VSS VDD
X0 net26 SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X1 net26 E VSS VSS LPNFET W=0.2U L=0.12U M=1 
X10 hnet28 cn net33 VDD LPPFET W=1U L=0.12U M=1 
X11 VDD net40 hnet28 VDD LPPFET W=1U L=0.12U M=1 
X12 hnet32 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X13 net33 cn hnet32 VSS LPNFET W=0.2U L=0.12U M=1 
X14 hnet34 c net33 VDD LPPFET W=0.28U L=0.12U M=1 
X15 VDD m hnet34 VDD LPPFET W=0.28U L=0.12U M=1 
X16 VDD net26 net40 VDD LPPFET W=0.38U L=0.12U M=1 
X17 net40 net26 VSS VSS LPNFET W=0.28U L=0.12U M=1 
X18 VDD c cn VDD LPPFET W=0.28U L=0.12U M=1 
X19 cn c VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 VDD SE hnet14 VDD LPPFET W=0.36U L=0.12U M=1 
X20 VDD CK c VDD LPPFET W=0.78U L=0.12U M=1 
X21 c CK VSS VSS LPNFET W=0.56U L=0.12U M=1 
X22 VDD net33 m VDD LPPFET W=0.28U L=0.12U M=1 
X23 m net33 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 hnet14 E net26 VDD LPPFET W=0.36U L=0.12U M=1 
X4 ECK c VSS VSS LPNFET W=0.38U L=0.12U M=1 
X5 ECK net33 VSS VSS LPNFET W=0.38U L=0.12U M=1 
X6 VDD c hnet20 VDD LPPFET W=1.3U L=0.12U M=1 
X7 hnet20 net33 ECK VDD LPPFET W=1.3U L=0.12U M=1 
X8 hnet26 net40 VSS VSS LPNFET W=0.72U L=0.12U M=1 
X9 net33 c hnet26 VSS LPNFET W=0.72U L=0.12U M=1 
.ENDS TLATNTSCAX2TS 

**** 
*.SUBCKT TLATNTSCAX3TS ECK CK E SE 
.SUBCKT TLATNTSCAX3TS ECK CK E SE VSS VDD
X0 net26 SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X1 net26 E VSS VSS LPNFET W=0.2U L=0.12U M=1 
X10 hnet25 net40 VSS VSS LPNFET W=0.84U L=0.12U M=1 
X11 net33 c hnet25 VSS LPNFET W=0.84U L=0.12U M=1 
X12 hnet27 cn net33 VDD LPPFET W=1.26U L=0.12U M=1 
X13 VDD net40 hnet27 VDD LPPFET W=1.26U L=0.12U M=1 
X14 hnet31 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X15 net33 cn hnet31 VSS LPNFET W=0.2U L=0.12U M=1 
X16 hnet33 c net33 VDD LPPFET W=0.28U L=0.12U M=1 
X17 VDD m hnet33 VDD LPPFET W=0.28U L=0.12U M=1 
X18 VDD net26 net40 VDD LPPFET W=0.5U L=0.12U M=1 
X19 net40 net26 VSS VSS LPNFET W=0.36U L=0.12U M=1 
X2 VDD SE hnet14 VDD LPPFET W=0.36U L=0.12U M=1 
X20 VDD c cn VDD LPPFET W=0.3U L=0.12U M=1 
X21 cn c VSS VSS LPNFET W=0.22U L=0.12U M=1 
X22 VDD CK c VDD LPPFET W=1U L=0.12U M=1 
X23 c CK VSS VSS LPNFET W=0.72U L=0.12U M=1 
X24 VDD net33 m VDD LPPFET W=0.28U L=0.12U M=1 
X25 m net33 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 hnet14 E net26 VDD LPPFET W=0.36U L=0.12U M=1 
X4 ECK c VSS VSS LPNFET W=0.56U L=0.12U M=1 
X5 ECK net33 VSS VSS LPNFET W=0.56U L=0.12U M=1 
X6 VDD c hnet21 VDD LPPFET W=0.96U L=0.12U M=1 
X7 hnet21 net33 ECK VDD LPPFET W=0.96U L=0.12U M=1 
X8 VDD c hnet19 VDD LPPFET W=0.96U L=0.12U M=1 
X9 hnet19 net33 ECK VDD LPPFET W=0.96U L=0.12U M=1 
.ENDS TLATNTSCAX3TS 

**** 
*.SUBCKT TLATNTSCAX4TS ECK CK E SE 
.SUBCKT TLATNTSCAX4TS ECK CK E SE VSS VDD
X0 net26 SE VSS VSS LPNFET W=0.2U L=0.12U M=1 
X1 net26 E VSS VSS LPNFET W=0.2U L=0.12U M=1 
X10 hnet25 net40 VSS VSS LPNFET W=0.64U L=0.12U M=1 
X11 hnet26 net40 VSS VSS LPNFET W=0.64U L=0.12U M=1 
X12 net33 c hnet25 VSS LPNFET W=0.64U L=0.12U M=1 
X13 net33 c hnet26 VSS LPNFET W=0.64U L=0.12U M=1 
X14 hnet31 cn net33 VDD LPPFET W=0.88U L=0.12U M=1 
X15 hnet29 cn net33 VDD LPPFET W=0.88U L=0.12U M=1 
X16 VDD net40 hnet31 VDD LPPFET W=0.88U L=0.12U M=1 
X17 VDD net40 hnet29 VDD LPPFET W=0.88U L=0.12U M=1 
X18 hnet33 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X19 net33 cn hnet33 VSS LPNFET W=0.2U L=0.12U M=1 
X2 VDD SE hnet14 VDD LPPFET W=0.36U L=0.12U M=1 
X20 hnet35 c net33 VDD LPPFET W=0.28U L=0.12U M=1 
X21 VDD m hnet35 VDD LPPFET W=0.28U L=0.12U M=1 
X22 VDD net26 net40 VDD LPPFET W=0.7U L=0.12U M=1 
X23 net40 net26 VSS VSS LPNFET W=0.5U L=0.12U M=1 
X24 VDD c cn VDD LPPFET W=0.42U L=0.12U M=1 
X25 cn c VSS VSS LPNFET W=0.3U L=0.12U M=1 
X26 VDD CK c VDD LPPFET W=1.36U L=0.12U M=1 
X27 c CK VSS VSS LPNFET W=0.92U L=0.12U M=1 
X28 VDD net33 m VDD LPPFET W=0.28U L=0.12U M=1 
X29 m net33 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 hnet14 E net26 VDD LPPFET W=0.36U L=0.12U M=1 
X4 ECK c VSS VSS LPNFET W=0.74U L=0.12U M=1 
X5 ECK net33 VSS VSS LPNFET W=0.74U L=0.12U M=1 
X6 VDD c hnet21 VDD LPPFET W=1.28U L=0.12U M=1 
X7 hnet21 net33 ECK VDD LPPFET W=1.28U L=0.12U M=1 
X8 VDD c hnet19 VDD LPPFET W=1.28U L=0.12U M=1 
X9 hnet19 net33 ECK VDD LPPFET W=1.28U L=0.12U M=1 
.ENDS TLATNTSCAX4TS 

**** 
*.SUBCKT TLATNTSCAX6TS ECK CK E SE 
.SUBCKT TLATNTSCAX6TS ECK CK E SE VSS VDD
X0 hnet15 net40 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X1 hnet17 net40 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X10 VDD net40 hnet18 VDD LPPFET W=0.84U L=0.12U M=1 
X11 VDD net40 hnet14 VDD LPPFET W=0.84U L=0.12U M=1 
X12 net30 SE VSS VSS LPNFET W=0.3U L=0.12U M=1 
X13 net30 E VSS VSS LPNFET W=0.3U L=0.12U M=1 
X14 VDD SE hnet26 VDD LPPFET W=0.54U L=0.12U M=1 
X15 hnet26 E net30 VDD LPPFET W=0.54U L=0.12U M=1 
X16 ECK c VSS VSS LPNFET W=1.12U L=0.12U M=1 
X17 ECK net27 VSS VSS LPNFET W=1.12U L=0.12U M=1 
X18 VDD c hnet31 VDD LPPFET W=1.28U L=0.12U M=1 
X19 hnet31 net27 ECK VDD LPPFET W=1.28U L=0.12U M=1 
X2 hnet22 net40 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X20 VDD c hnet29 VDD LPPFET W=1.28U L=0.12U M=1 
X21 hnet29 net27 ECK VDD LPPFET W=1.28U L=0.12U M=1 
X22 VDD c hnet32 VDD LPPFET W=1.28U L=0.12U M=1 
X23 hnet32 net27 ECK VDD LPPFET W=1.28U L=0.12U M=1 
X24 hnet36 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X25 net27 cn hnet36 VSS LPNFET W=0.2U L=0.12U M=1 
X26 hnet38 c net27 VDD LPPFET W=0.28U L=0.12U M=1 
X27 VDD m hnet38 VDD LPPFET W=0.28U L=0.12U M=1 
X28 VDD net30 net40 VDD LPPFET W=1.02U L=0.12U M=1 
X29 net40 net30 VSS VSS LPNFET W=0.74U L=0.12U M=1 
X3 net27 c hnet15 VSS LPNFET W=0.6U L=0.12U M=1 
X30 VDD c cn VDD LPPFET W=0.56U L=0.12U M=1 
X31 cn c VSS VSS LPNFET W=0.4U L=0.12U M=1 
X32 VDD CK c VDD LPPFET W=1.92U L=0.12U M=1 
X33 c CK VSS VSS LPNFET W=1.38U L=0.12U M=1 
X34 VDD net27 m VDD LPPFET W=0.28U L=0.12U M=1 
X35 m net27 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X4 net27 c hnet17 VSS LPNFET W=0.6U L=0.12U M=1 
X5 net27 c hnet22 VSS LPNFET W=0.6U L=0.12U M=1 
X6 hnet16 cn net27 VDD LPPFET W=0.84U L=0.12U M=1 
X7 hnet18 cn net27 VDD LPPFET W=0.84U L=0.12U M=1 
X8 hnet14 cn net27 VDD LPPFET W=0.84U L=0.12U M=1 
X9 VDD net40 hnet16 VDD LPPFET W=0.84U L=0.12U M=1 
.ENDS TLATNTSCAX6TS 

**** 
*.SUBCKT TLATNTSCAX8TS ECK CK E SE 
.SUBCKT TLATNTSCAX8TS ECK CK E SE VSS VDD
X0 ECK c VSS VSS LPNFET W=1.84U L=0.12U M=1 
X1 ECK net49 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X10 VDD c hnet20 VDD LPPFET W=1.3U L=0.12U M=1 
X11 hnet20 net49 ECK VDD LPPFET W=1.3U L=0.12U M=1 
X12 VDD c hnet17 VDD LPPFET W=1.3U L=0.12U M=1 
X13 hnet17 net49 ECK VDD LPPFET W=1.3U L=0.12U M=1 
X14 VDD c hnet25 VDD LPPFET W=1.3U L=0.12U M=1 
X15 hnet25 net49 ECK VDD LPPFET W=1.3U L=0.12U M=1 
X16 net49 c net37 VSS LPNFET W=0.92U L=0.12U M=1 
X17 net37 net59 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X18 VDD net59 net47 VDD LPPFET W=1.12U L=0.12U M=1 
X19 net47 cn net49 VDD LPPFET W=1.12U L=0.12U M=1 
X2 VDD c hnet23 VDD LPPFET W=1.3U L=0.12U M=1 
X20 hnet28 net59 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X21 hnet30 net59 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X22 hnet37 net59 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X23 hnet29 net59 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X24 net49 c hnet28 VSS LPNFET W=0.6U L=0.12U M=1 
X25 net49 c hnet30 VSS LPNFET W=0.6U L=0.12U M=1 
X26 net49 c hnet37 VSS LPNFET W=0.6U L=0.12U M=1 
X27 net49 c hnet29 VSS LPNFET W=0.6U L=0.12U M=1 
X28 hnet35 cn net49 VDD LPPFET W=0.86U L=0.12U M=1 
X29 hnet38 cn net49 VDD LPPFET W=0.86U L=0.12U M=1 
X3 hnet23 net49 ECK VDD LPPFET W=1.3U L=0.12U M=1 
X30 hnet31 cn net49 VDD LPPFET W=0.86U L=0.12U M=1 
X31 hnet36 cn net49 VDD LPPFET W=0.86U L=0.12U M=1 
X32 VDD net59 hnet35 VDD LPPFET W=0.86U L=0.12U M=1 
X33 VDD net59 hnet38 VDD LPPFET W=0.86U L=0.12U M=1 
X34 VDD net59 hnet31 VDD LPPFET W=0.86U L=0.12U M=1 
X35 VDD net59 hnet36 VDD LPPFET W=0.86U L=0.12U M=1 
X36 net52 SE VSS VSS LPNFET W=0.6U L=0.12U M=1 
X37 net52 E VSS VSS LPNFET W=0.6U L=0.12U M=1 
X38 VDD SE hnet40 VDD LPPFET W=1.1U L=0.12U M=1 
X39 hnet40 E net52 VDD LPPFET W=1.1U L=0.12U M=1 
X4 VDD c hnet18 VDD LPPFET W=1.3U L=0.12U M=1 
X40 hnet44 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X41 net49 cn hnet44 VSS LPNFET W=0.2U L=0.12U M=1 
X42 hnet46 c net49 VDD LPPFET W=0.28U L=0.12U M=1 
X43 VDD m hnet46 VDD LPPFET W=0.28U L=0.12U M=1 
X44 VDD net52 net59 VDD LPPFET W=2.06U L=0.12U M=1 
X45 net59 net52 VSS VSS LPNFET W=1.48U L=0.12U M=1 
X46 VDD c cn VDD LPPFET W=1.08U L=0.12U M=1 
X47 cn c VSS VSS LPNFET W=0.74U L=0.12U M=1 
X48 VDD CK c VDD LPPFET W=3.9U L=0.12U M=1 
X49 c CK VSS VSS LPNFET W=2.76U L=0.12U M=1 
X5 hnet18 net49 ECK VDD LPPFET W=1.3U L=0.12U M=1 
X50 VDD net49 m VDD LPPFET W=0.28U L=0.12U M=1 
X51 m net49 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X6 VDD c hnet22 VDD LPPFET W=1.3U L=0.12U M=1 
X7 hnet22 net49 ECK VDD LPPFET W=1.3U L=0.12U M=1 
X8 VDD c hnet21 VDD LPPFET W=1.3U L=0.12U M=1 
X9 hnet21 net49 ECK VDD LPPFET W=1.3U L=0.12U M=1 
.ENDS TLATNTSCAX8TS 

**** 
*.SUBCKT TLATNX1TS Q QN D GN 
.SUBCKT TLATNX1TS Q QN D GN VSS VDD
X0 hnet12 D VSS VSS LPNFET W=0.48U L=0.12U M=1 
X1 nmin c hnet12 VSS LPNFET W=0.48U L=0.12U M=1 
X10 VDD GN c VDD LPPFET W=0.34U L=0.12U M=1 
X11 c GN VSS VSS LPNFET W=0.28U L=0.12U M=1 
X12 VDD nmin Q VDD LPPFET W=0.64U L=0.12U M=1 
X13 Q nmin VSS VSS LPNFET W=0.44U L=0.12U M=1 
X14 VDD m QN VDD LPPFET W=0.64U L=0.12U M=1 
X15 QN m VSS VSS LPNFET W=0.46U L=0.12U M=1 
X16 VDD nmin m VDD LPPFET W=0.28U L=0.12U M=1 
X17 m nmin VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 hnet14 cn nmin VDD LPPFET W=0.72U L=0.12U M=1 
X3 VDD D hnet14 VDD LPPFET W=0.72U L=0.12U M=1 
X4 hnet20 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X5 nmin cn hnet20 VSS LPNFET W=0.2U L=0.12U M=1 
X6 hnet22 c nmin VDD LPPFET W=0.28U L=0.12U M=1 
X7 VDD m hnet22 VDD LPPFET W=0.28U L=0.12U M=1 
X8 VDD c cn VDD LPPFET W=0.28U L=0.12U M=1 
X9 cn c VSS VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS TLATNX1TS 

**** 
*.SUBCKT TLATNX2TS Q QN D GN 
.SUBCKT TLATNX2TS Q QN D GN VSS VDD
X0 hnet12 D VSS VSS LPNFET W=0.84U L=0.12U M=1 
X1 nmin c hnet12 VSS LPNFET W=0.84U L=0.12U M=1 
X10 VDD GN c VDD LPPFET W=0.42U L=0.12U M=1 
X11 c GN VSS VSS LPNFET W=0.3U L=0.12U M=1 
X12 VDD nmin Q VDD LPPFET W=1.28U L=0.12U M=1 
X13 Q nmin VSS VSS LPNFET W=0.92U L=0.12U M=1 
X14 VDD m QN VDD LPPFET W=1.28U L=0.12U M=1 
X15 QN m VSS VSS LPNFET W=0.92U L=0.12U M=1 
X16 VDD nmin m VDD LPPFET W=0.44U L=0.12U M=1 
X17 m nmin VSS VSS LPNFET W=0.32U L=0.12U M=1 
X2 hnet14 cn nmin VDD LPPFET W=1.26U L=0.12U M=1 
X3 VDD D hnet14 VDD LPPFET W=1.26U L=0.12U M=1 
X4 hnet20 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X5 nmin cn hnet20 VSS LPNFET W=0.2U L=0.12U M=1 
X6 hnet22 c nmin VDD LPPFET W=0.28U L=0.12U M=1 
X7 VDD m hnet22 VDD LPPFET W=0.28U L=0.12U M=1 
X8 VDD c cn VDD LPPFET W=0.3U L=0.12U M=1 
X9 cn c VSS VSS LPNFET W=0.22U L=0.12U M=1 
.ENDS TLATNX2TS 

**** 
*.SUBCKT TLATNX4TS Q QN D GN 
.SUBCKT TLATNX4TS Q QN D GN VSS VDD
X0 hnet12 D VSS VSS LPNFET W=0.92U L=0.12U M=1 
X1 hnet13 D VSS VSS LPNFET W=0.92U L=0.12U M=1 
X10 hnet24 c nmin VDD LPPFET W=0.28U L=0.12U M=1 
X11 VDD m hnet24 VDD LPPFET W=0.28U L=0.12U M=1 
X12 VDD c cn VDD LPPFET W=0.56U L=0.12U M=1 
X13 cn c VSS VSS LPNFET W=0.4U L=0.12U M=1 
X14 VDD GN c VDD LPPFET W=0.78U L=0.12U M=1 
X15 c GN VSS VSS LPNFET W=0.56U L=0.12U M=1 
X16 VDD nmin Q VDD LPPFET W=2.48U L=0.12U M=1 
X17 Q nmin VSS VSS LPNFET W=1.84U L=0.12U M=1 
X18 VDD m QN VDD LPPFET W=2.48U L=0.12U M=1 
X19 QN m VSS VSS LPNFET W=1.84U L=0.12U M=1 
X2 nmin c hnet12 VSS LPNFET W=0.92U L=0.12U M=1 
X20 VDD nmin m VDD LPPFET W=0.8U L=0.12U M=1 
X21 m nmin VSS VSS LPNFET W=0.58U L=0.12U M=1 
X3 nmin c hnet13 VSS LPNFET W=0.92U L=0.12U M=1 
X4 hnet20 cn nmin VDD LPPFET W=1.2U L=0.12U M=1 
X5 hnet17 cn nmin VDD LPPFET W=1.2U L=0.12U M=1 
X6 VDD D hnet20 VDD LPPFET W=1.2U L=0.12U M=1 
X7 VDD D hnet17 VDD LPPFET W=1.2U L=0.12U M=1 
X8 hnet22 m VSS VSS LPNFET W=0.18U L=0.12U M=1 
X9 nmin cn hnet22 VSS LPNFET W=0.18U L=0.12U M=1 
.ENDS TLATNX4TS 

**** 
*.SUBCKT TLATNXLTS Q QN D GN 
.SUBCKT TLATNXLTS Q QN D GN VSS VDD
X0 hnet12 D VSS VSS LPNFET W=0.2U L=0.12U M=1 
X1 nmin c hnet12 VSS LPNFET W=0.2U L=0.12U M=1 
X10 VDD GN c VDD LPPFET W=0.28U L=0.12U M=1 
X11 c GN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X12 VDD nmin Q VDD LPPFET W=0.42U L=0.12U M=1 
X13 Q nmin VSS VSS LPNFET W=0.24U L=0.12U M=1 
X14 VDD m QN VDD LPPFET W=0.42U L=0.12U M=1 
X15 QN m VSS VSS LPNFET W=0.24U L=0.12U M=1 
X16 VDD nmin m VDD LPPFET W=0.28U L=0.12U M=1 
X17 m nmin VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 hnet14 cn nmin VDD LPPFET W=0.28U L=0.12U M=1 
X3 VDD D hnet14 VDD LPPFET W=0.28U L=0.12U M=1 
X4 hnet20 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X5 nmin cn hnet20 VSS LPNFET W=0.2U L=0.12U M=1 
X6 hnet22 c nmin VDD LPPFET W=0.28U L=0.12U M=1 
X7 VDD m hnet22 VDD LPPFET W=0.28U L=0.12U M=1 
X8 VDD c cn VDD LPPFET W=0.28U L=0.12U M=1 
X9 cn c VSS VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS TLATNXLTS 

**** 
*.SUBCKT TLATSRX1TS Q QN D G RN SN 
.SUBCKT TLATSRX1TS Q QN D G RN SN VSS VDD
X0 VDD D hnet20 VDD LPPFET W=0.6U L=0.12U M=1 
X1 hnet20 nms hnet25 VDD LPPFET W=0.6U L=0.12U M=1 
X10 VDD pm Q VDD LPPFET W=0.56U L=0.12U M=1 
X11 Q pm VSS VSS LPNFET W=0.42U L=0.12U M=1 
X12 VDD SN nms VDD LPPFET W=0.42U L=0.12U M=1 
X13 nms SN VSS VSS LPNFET W=0.3U L=0.12U M=1 
X14 VDD cn c VDD LPPFET W=0.26U L=0.12U M=1 
X15 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X16 VDD G cn VDD LPPFET W=0.38U L=0.12U M=1 
X17 cn G VSS VSS LPNFET W=0.28U L=0.12U M=1 
X18 VDD pm m VDD LPPFET W=0.3U L=0.12U M=1 
X19 m pm VSS VSS LPNFET W=0.22U L=0.12U M=1 
X2 hnet25 cn pm VDD LPPFET W=0.6U L=0.12U M=1 
X20 net65 nms net71 VDD LPPFET W=0.36U L=0.12U M=1 
X21 pm c net65 VDD LPPFET W=0.36U L=0.12U M=1 
X22 net71 m VDD VDD LPPFET W=0.36U L=0.12U M=1 
X23 net74 RN net77 VSS LPNFET W=0.32U L=0.12U M=1 
X24 net77 m VSS VSS LPNFET W=0.32U L=0.12U M=1 
X25 pm cn net74 VSS LPNFET W=0.32U L=0.12U M=1 
X26 pm nms VSS VSS LPNFET W=0.28U L=0.12U M=1 
X3 hnet31 D VSS VSS LPNFET W=0.42U L=0.12U M=1 
X4 hnet26 RN hnet31 VSS LPNFET W=0.42U L=0.12U M=1 
X5 pm c hnet26 VSS LPNFET W=0.42U L=0.12U M=1 
X6 VDD RN hnet35 VDD LPPFET W=0.5U L=0.12U M=1 
X7 hnet35 nms pm VDD LPPFET W=0.5U L=0.12U M=1 
X8 VDD m QN VDD LPPFET W=0.56U L=0.12U M=1 
X9 QN m VSS VSS LPNFET W=0.46U L=0.12U M=1 
.ENDS TLATSRX1TS 

**** 
*.SUBCKT TLATSRX2TS Q QN D G RN SN 
.SUBCKT TLATSRX2TS Q QN D G RN SN VSS VDD
X0 VDD D hnet20 VDD LPPFET W=1.12U L=0.12U M=1 
X1 hnet20 nms hnet25 VDD LPPFET W=1.12U L=0.12U M=1 
X10 VDD pm Q VDD LPPFET W=1.28U L=0.12U M=1 
X11 Q pm VSS VSS LPNFET W=0.9U L=0.12U M=1 
X12 VDD SN nms VDD LPPFET W=0.66U L=0.12U M=1 
X13 nms SN VSS VSS LPNFET W=0.48U L=0.12U M=1 
X14 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X15 c cn VSS VSS LPNFET W=0.22U L=0.12U M=1 
X16 VDD G cn VDD LPPFET W=0.42U L=0.12U M=1 
X17 cn G VSS VSS LPNFET W=0.28U L=0.12U M=1 
X18 VDD pm m VDD LPPFET W=0.48U L=0.12U M=1 
X19 m pm VSS VSS LPNFET W=0.34U L=0.12U M=1 
X2 hnet25 cn pm VDD LPPFET W=1.12U L=0.12U M=1 
X20 net65 nms net71 VDD LPPFET W=0.36U L=0.12U M=1 
X21 pm c net65 VDD LPPFET W=0.36U L=0.12U M=1 
X22 net71 m VDD VDD LPPFET W=0.36U L=0.12U M=1 
X23 net74 RN net77 VSS LPNFET W=0.32U L=0.12U M=1 
X24 net77 m VSS VSS LPNFET W=0.32U L=0.12U M=1 
X25 pm cn net74 VSS LPNFET W=0.32U L=0.12U M=1 
X26 pm nms VSS VSS LPNFET W=0.5U L=0.12U M=1 
X3 hnet31 D VSS VSS LPNFET W=0.64U L=0.12U M=1 
X4 hnet26 RN hnet31 VSS LPNFET W=0.64U L=0.12U M=1 
X5 pm c hnet26 VSS LPNFET W=0.64U L=0.12U M=1 
X6 VDD RN hnet35 VDD LPPFET W=0.88U L=0.12U M=1 
X7 hnet35 nms pm VDD LPPFET W=0.88U L=0.12U M=1 
X8 VDD m QN VDD LPPFET W=1.28U L=0.12U M=1 
X9 QN m VSS VSS LPNFET W=0.9U L=0.12U M=1 
.ENDS TLATSRX2TS 

**** 
*.SUBCKT TLATSRX4TS Q QN D G RN SN 
.SUBCKT TLATSRX4TS Q QN D G RN SN VSS VDD
X0 VDD D hnet21 VDD LPPFET W=0.98U L=0.12U M=1 
X1 hnet21 nms hnet20 VDD LPPFET W=0.98U L=0.12U M=1 
X10 hnet36 RN hnet37 VSS LPNFET W=0.48U L=0.12U M=1 
X11 pm c hnet36 VSS LPNFET W=0.48U L=0.12U M=1 
X12 hnet31 D VSS VSS LPNFET W=0.48U L=0.12U M=1 
X13 hnet29 RN hnet31 VSS LPNFET W=0.48U L=0.12U M=1 
X14 pm c hnet29 VSS LPNFET W=0.48U L=0.12U M=1 
X15 VDD RN hnet42 VDD LPPFET W=0.92U L=0.12U M=1 
X16 hnet42 nms pm VDD LPPFET W=0.92U L=0.12U M=1 
X17 VDD RN hnet39 VDD LPPFET W=0.92U L=0.12U M=1 
X18 hnet39 nms pm VDD LPPFET W=0.92U L=0.12U M=1 
X19 VDD m QN VDD LPPFET W=2.56U L=0.12U M=1 
X2 hnet20 cn pm VDD LPPFET W=0.98U L=0.12U M=1 
X20 QN m VSS VSS LPNFET W=1.84U L=0.12U M=1 
X21 VDD pm Q VDD LPPFET W=2.56U L=0.12U M=1 
X22 Q pm VSS VSS LPNFET W=1.84U L=0.12U M=1 
X23 VDD SN nms VDD LPPFET W=1.22U L=0.12U M=1 
X24 nms SN VSS VSS LPNFET W=0.88U L=0.12U M=1 
X25 VDD cn c VDD LPPFET W=0.5U L=0.12U M=1 
X26 c cn VSS VSS LPNFET W=0.36U L=0.12U M=1 
X27 VDD G cn VDD LPPFET W=0.7U L=0.12U M=1 
X28 cn G VSS VSS LPNFET W=0.5U L=0.12U M=1 
X29 VDD pm m VDD LPPFET W=0.84U L=0.12U M=1 
X3 VDD D hnet23 VDD LPPFET W=0.98U L=0.12U M=1 
X30 m pm VSS VSS LPNFET W=0.6U L=0.12U M=1 
X31 net65 nms net71 VDD LPPFET W=0.32U L=0.12U M=1 
X32 pm c net65 VDD LPPFET W=0.32U L=0.12U M=1 
X33 net71 m VDD VDD LPPFET W=0.32U L=0.12U M=1 
X34 net74 RN net77 VSS LPNFET W=0.32U L=0.12U M=1 
X35 net77 m VSS VSS LPNFET W=0.32U L=0.12U M=1 
X36 pm cn net74 VSS LPNFET W=0.32U L=0.12U M=1 
X37 pm nms VSS VSS LPNFET W=0.92U L=0.12U M=1 
X4 hnet23 nms hnet24 VDD LPPFET W=0.98U L=0.12U M=1 
X5 hnet24 cn pm VDD LPPFET W=0.98U L=0.12U M=1 
X6 hnet35 D VSS VSS LPNFET W=0.48U L=0.12U M=1 
X7 hnet28 RN hnet35 VSS LPNFET W=0.48U L=0.12U M=1 
X8 pm c hnet28 VSS LPNFET W=0.48U L=0.12U M=1 
X9 hnet37 D VSS VSS LPNFET W=0.48U L=0.12U M=1 
.ENDS TLATSRX4TS 

**** 
*.SUBCKT TLATSRXLTS Q QN D G RN SN 
.SUBCKT TLATSRXLTS Q QN D G RN SN VSS VDD
X0 VDD D hnet20 VDD LPPFET W=0.36U L=0.12U M=1 
X1 hnet20 nms hnet25 VDD LPPFET W=0.36U L=0.12U M=1 
X10 VDD pm Q VDD LPPFET W=0.42U L=0.12U M=1 
X11 Q pm VSS VSS LPNFET W=0.24U L=0.12U M=1 
X12 VDD SN nms VDD LPPFET W=0.28U L=0.12U M=1 
X13 nms SN VSS VSS LPNFET W=0.2U L=0.12U M=1 
X14 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X15 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
X16 VDD G cn VDD LPPFET W=0.28U L=0.12U M=1 
X17 cn G VSS VSS LPNFET W=0.2U L=0.12U M=1 
X18 VDD pm m VDD LPPFET W=0.28U L=0.12U M=1 
X19 m pm VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 hnet25 cn pm VDD LPPFET W=0.36U L=0.12U M=1 
X20 net65 nms net71 VDD LPPFET W=0.36U L=0.12U M=1 
X21 pm c net65 VDD LPPFET W=0.36U L=0.12U M=1 
X22 net71 m VDD VDD LPPFET W=0.36U L=0.12U M=1 
X23 net74 RN net77 VSS LPNFET W=0.32U L=0.12U M=1 
X24 net77 m VSS VSS LPNFET W=0.32U L=0.12U M=1 
X25 pm cn net74 VSS LPNFET W=0.32U L=0.12U M=1 
X26 pm nms VSS VSS LPNFET W=0.2U L=0.12U M=1 
X3 hnet31 D VSS VSS LPNFET W=0.32U L=0.12U M=1 
X4 hnet26 RN hnet31 VSS LPNFET W=0.32U L=0.12U M=1 
X5 pm c hnet26 VSS LPNFET W=0.32U L=0.12U M=1 
X6 VDD RN hnet35 VDD LPPFET W=0.3U L=0.12U M=1 
X7 hnet35 nms pm VDD LPPFET W=0.3U L=0.12U M=1 
X8 VDD m QN VDD LPPFET W=0.42U L=0.12U M=1 
X9 QN m VSS VSS LPNFET W=0.24U L=0.12U M=1 
.ENDS TLATSRXLTS 

**** 
*.SUBCKT TLATX1TS Q QN D G 
.SUBCKT TLATX1TS Q QN D G VSS VDD
X0 hnet12 D VSS VSS LPNFET W=0.48U L=0.12U M=1 
X1 pm c hnet12 VSS LPNFET W=0.48U L=0.12U M=1 
X10 VDD G cn VDD LPPFET W=0.38U L=0.12U M=1 
X11 cn G VSS VSS LPNFET W=0.28U L=0.12U M=1 
X12 VDD pm Q VDD LPPFET W=0.64U L=0.12U M=1 
X13 Q pm VSS VSS LPNFET W=0.46U L=0.12U M=1 
X14 VDD m QN VDD LPPFET W=0.64U L=0.12U M=1 
X15 QN m VSS VSS LPNFET W=0.46U L=0.12U M=1 
X16 VDD pm m VDD LPPFET W=0.28U L=0.12U M=1 
X17 m pm VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 hnet14 cn pm VDD LPPFET W=0.72U L=0.12U M=1 
X3 VDD D hnet14 VDD LPPFET W=0.72U L=0.12U M=1 
X4 hnet20 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X5 pm cn hnet20 VSS LPNFET W=0.2U L=0.12U M=1 
X6 hnet22 c pm VDD LPPFET W=0.28U L=0.12U M=1 
X7 VDD m hnet22 VDD LPPFET W=0.28U L=0.12U M=1 
X8 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X9 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS TLATX1TS 

**** 
*.SUBCKT TLATX2TS Q QN D G 
.SUBCKT TLATX2TS Q QN D G VSS VDD
X0 hnet12 D VSS VSS LPNFET W=0.84U L=0.12U M=1 
X1 pm c hnet12 VSS LPNFET W=0.84U L=0.12U M=1 
X10 VDD G cn VDD LPPFET W=0.42U L=0.12U M=1 
X11 cn G VSS VSS LPNFET W=0.3U L=0.12U M=1 
X12 VDD pm Q VDD LPPFET W=1.28U L=0.12U M=1 
X13 Q pm VSS VSS LPNFET W=0.92U L=0.12U M=1 
X14 VDD m QN VDD LPPFET W=1.28U L=0.12U M=1 
X15 QN m VSS VSS LPNFET W=0.92U L=0.12U M=1 
X16 VDD pm m VDD LPPFET W=0.44U L=0.12U M=1 
X17 m pm VSS VSS LPNFET W=0.32U L=0.12U M=1 
X2 hnet14 cn pm VDD LPPFET W=1.26U L=0.12U M=1 
X3 VDD D hnet14 VDD LPPFET W=1.26U L=0.12U M=1 
X4 hnet20 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X5 pm cn hnet20 VSS LPNFET W=0.2U L=0.12U M=1 
X6 hnet22 c pm VDD LPPFET W=0.28U L=0.12U M=1 
X7 VDD m hnet22 VDD LPPFET W=0.28U L=0.12U M=1 
X8 VDD cn c VDD LPPFET W=0.3U L=0.12U M=1 
X9 c cn VSS VSS LPNFET W=0.22U L=0.12U M=1 
.ENDS TLATX2TS 

**** 
*.SUBCKT TLATX4TS Q QN D G 
.SUBCKT TLATX4TS Q QN D G VSS VDD
X0 hnet12 D VSS VSS LPNFET W=0.66U L=0.12U M=1 
X1 hnet13 D VSS VSS LPNFET W=0.66U L=0.12U M=1 
X10 hnet24 c pm VDD LPPFET W=0.28U L=0.12U M=1 
X11 VDD m hnet24 VDD LPPFET W=0.28U L=0.12U M=1 
X12 VDD cn c VDD LPPFET W=0.56U L=0.12U M=1 
X13 c cn VSS VSS LPNFET W=0.4U L=0.12U M=1 
X14 VDD G cn VDD LPPFET W=0.78U L=0.12U M=1 
X15 cn G VSS VSS LPNFET W=0.56U L=0.12U M=1 
X16 VDD pm Q VDD LPPFET W=2.48U L=0.12U M=1 
X17 Q pm VSS VSS LPNFET W=1.84U L=0.12U M=1 
X18 VDD m QN VDD LPPFET W=2.48U L=0.12U M=1 
X19 QN m VSS VSS LPNFET W=1.84U L=0.12U M=1 
X2 pm c hnet12 VSS LPNFET W=0.66U L=0.12U M=1 
X20 VDD pm m VDD LPPFET W=0.8U L=0.12U M=1 
X21 m pm VSS VSS LPNFET W=0.52U L=0.12U M=1 
X3 pm c hnet13 VSS LPNFET W=0.66U L=0.12U M=1 
X4 hnet20 cn pm VDD LPPFET W=1.14U L=0.12U M=1 
X5 hnet17 cn pm VDD LPPFET W=1.14U L=0.12U M=1 
X6 VDD D hnet20 VDD LPPFET W=1.14U L=0.12U M=1 
X7 VDD D hnet17 VDD LPPFET W=1.14U L=0.12U M=1 
X8 hnet22 m VSS VSS LPNFET W=0.18U L=0.12U M=1 
X9 pm cn hnet22 VSS LPNFET W=0.18U L=0.12U M=1 
.ENDS TLATX4TS 

**** 
*.SUBCKT TLATXLTS Q QN D G 
.SUBCKT TLATXLTS Q QN D G VSS VDD
X0 hnet12 D VSS VSS LPNFET W=0.2U L=0.12U M=1 
X1 pm c hnet12 VSS LPNFET W=0.2U L=0.12U M=1 
X10 VDD G cn VDD LPPFET W=0.28U L=0.12U M=1 
X11 cn G VSS VSS LPNFET W=0.2U L=0.12U M=1 
X12 VDD pm Q VDD LPPFET W=0.42U L=0.12U M=1 
X13 Q pm VSS VSS LPNFET W=0.24U L=0.12U M=1 
X14 VDD m QN VDD LPPFET W=0.42U L=0.12U M=1 
X15 QN m VSS VSS LPNFET W=0.24U L=0.12U M=1 
X16 VDD pm m VDD LPPFET W=0.28U L=0.12U M=1 
X17 m pm VSS VSS LPNFET W=0.2U L=0.12U M=1 
X2 hnet14 cn pm VDD LPPFET W=0.28U L=0.12U M=1 
X3 VDD D hnet14 VDD LPPFET W=0.28U L=0.12U M=1 
X4 hnet20 m VSS VSS LPNFET W=0.2U L=0.12U M=1 
X5 pm cn hnet20 VSS LPNFET W=0.2U L=0.12U M=1 
X6 hnet22 c pm VDD LPPFET W=0.28U L=0.12U M=1 
X7 VDD m hnet22 VDD LPPFET W=0.28U L=0.12U M=1 
X8 VDD cn c VDD LPPFET W=0.28U L=0.12U M=1 
X9 c cn VSS VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS TLATXLTS 

**** 
*.SUBCKT XNOR2X1TS Y A B 
.SUBCKT XNOR2X1TS Y A B VSS VDD
X0 Y nmin1 net35 VDD LPPFET W=0.78U L=0.12U M=1 
X1 Y A nmin2 VDD LPPFET W=0.78U L=0.12U M=1 
X2 Y A net35 VSS LPNFET W=0.56U L=0.12U M=1 
X3 Y nmin1 nmin2 VSS LPNFET W=0.56U L=0.12U M=1 
X4 VDD A nmin1 VDD LPPFET W=0.3U L=0.12U M=1 
X5 nmin1 A VSS VSS LPNFET W=0.22U L=0.12U M=1 
X6 VDD nmin2 net35 VDD LPPFET W=0.78U L=0.12U M=1 
X7 net35 nmin2 VSS VSS LPNFET W=0.56U L=0.12U M=1 
X8 VDD B nmin2 VDD LPPFET W=0.72U L=0.12U M=1 
X9 nmin2 B VSS VSS LPNFET W=0.56U L=0.12U M=1 
.ENDS XNOR2X1TS 

**** 
*.SUBCKT XNOR2X2TS Y A B 
.SUBCKT XNOR2X2TS Y A B VSS VDD
X0 Y nmin1 net35 VDD LPPFET W=1.56U L=0.12U M=1 
X1 Y A nmin2 VDD LPPFET W=1.56U L=0.12U M=1 
X2 Y A net35 VSS LPNFET W=1.1U L=0.12U M=1 
X3 Y nmin1 nmin2 VSS LPNFET W=1.1U L=0.12U M=1 
X4 VDD A nmin1 VDD LPPFET W=0.62U L=0.12U M=1 
X5 nmin1 A VSS VSS LPNFET W=0.44U L=0.12U M=1 
X6 VDD nmin2 net35 VDD LPPFET W=1.56U L=0.12U M=1 
X7 net35 nmin2 VSS VSS LPNFET W=1.1U L=0.12U M=1 
X8 VDD B nmin2 VDD LPPFET W=1.56U L=0.12U M=1 
X9 nmin2 B VSS VSS LPNFET W=1.1U L=0.12U M=1 
.ENDS XNOR2X2TS 

**** 
*.SUBCKT XNOR2X4TS Y A B 
.SUBCKT XNOR2X4TS Y A B VSS VDD
X0 Y nmin1 net35 VDD LPPFET W=3.12U L=0.12U M=1 
X1 Y A nmin2 VDD LPPFET W=3.12U L=0.12U M=1 
X2 Y A net35 VSS LPNFET W=2.1U L=0.12U M=1 
X3 Y nmin1 nmin2 VSS LPNFET W=2.1U L=0.12U M=1 
X4 VDD A nmin1 VDD LPPFET W=1.22U L=0.12U M=1 
X5 nmin1 A VSS VSS LPNFET W=0.88U L=0.12U M=1 
X6 VDD nmin2 net35 VDD LPPFET W=3.12U L=0.12U M=1 
X7 net35 nmin2 VSS VSS LPNFET W=2.1U L=0.12U M=1 
X8 VDD B nmin2 VDD LPPFET W=3.12U L=0.12U M=1 
X9 nmin2 B VSS VSS LPNFET W=2.16U L=0.12U M=1 
.ENDS XNOR2X4TS 

**** 
*.SUBCKT XNOR2XLTS Y A B 
.SUBCKT XNOR2XLTS Y A B VSS VDD
X0 Y nmin1 net35 VDD LPPFET W=0.4U L=0.12U M=1 
X1 Y A nmin2 VDD LPPFET W=0.4U L=0.12U M=1 
X2 Y A net35 VSS LPNFET W=0.28U L=0.12U M=1 
X3 Y nmin1 nmin2 VSS LPNFET W=0.28U L=0.12U M=1 
X4 VDD A nmin1 VDD LPPFET W=0.28U L=0.12U M=1 
X5 nmin1 A VSS VSS LPNFET W=0.2U L=0.12U M=1 
X6 VDD nmin2 net35 VDD LPPFET W=0.4U L=0.12U M=1 
X7 net35 nmin2 VSS VSS LPNFET W=0.28U L=0.12U M=1 
X8 VDD B nmin2 VDD LPPFET W=0.4U L=0.12U M=1 
X9 nmin2 B VSS VSS LPNFET W=0.28U L=0.12U M=1 
.ENDS XNOR2XLTS 

**** 
*.SUBCKT XNOR3X1TS Y A B C 
.SUBCKT XNOR3X1TS Y A B C VSS VDD
X0 VDD nmin1 net54 VDD LPPFET W=0.5U L=0.12U M=1 
X1 net54 nmin1 VSS VSS LPNFET W=0.36U L=0.12U M=1 
X10 net87 nmin2 nmin1 VDD LPPFET W=0.72U L=0.12U M=1 
X11 net87 B net54 VDD LPPFET W=0.5U L=0.12U M=1 
X12 net93 nmin3 net99 VDD LPPFET W=0.5U L=0.12U M=1 
X13 net93 C net87 VDD LPPFET W=0.5U L=0.12U M=1 
X14 net99 B nmin1 VDD LPPFET W=0.72U L=0.12U M=1 
X15 net99 nmin2 net54 VDD LPPFET W=0.5U L=0.12U M=1 
X16 net87 B nmin1 VSS LPNFET W=0.52U L=0.12U M=1 
X17 net87 nmin2 net54 VSS LPNFET W=0.36U L=0.12U M=1 
X18 net93 C net99 VSS LPNFET W=0.36U L=0.12U M=1 
X19 net93 nmin3 net87 VSS LPNFET W=0.36U L=0.12U M=1 
X2 VDD net93 Y VDD LPPFET W=0.64U L=0.12U M=1 
X20 net99 nmin2 nmin1 VSS LPNFET W=0.52U L=0.12U M=1 
X21 net99 B net54 VSS LPNFET W=0.36U L=0.12U M=1 
X3 Y net93 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X4 VDD C nmin3 VDD LPPFET W=0.28U L=0.12U M=1 
X5 nmin3 C VSS VSS LPNFET W=0.2U L=0.12U M=1 
X6 VDD B nmin2 VDD LPPFET W=0.5U L=0.12U M=1 
X7 nmin2 B VSS VSS LPNFET W=0.36U L=0.12U M=1 
X8 VDD A nmin1 VDD LPPFET W=0.72U L=0.12U M=1 
X9 nmin1 A VSS VSS LPNFET W=0.52U L=0.12U M=1 
.ENDS XNOR3X1TS 

**** 
*.SUBCKT XNOR3X2TS Y A B C 
.SUBCKT XNOR3X2TS Y A B C VSS VDD
X0 VDD nmin1 net54 VDD LPPFET W=0.96U L=0.12U M=1 
X1 net54 nmin1 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X10 net87 nmin2 nmin1 VDD LPPFET W=1.28U L=0.12U M=1 
X11 net87 B net54 VDD LPPFET W=1.02U L=0.12U M=1 
X12 net93 nmin3 net99 VDD LPPFET W=0.98U L=0.12U M=1 
X13 net93 C net87 VDD LPPFET W=1.02U L=0.12U M=1 
X14 net99 B nmin1 VDD LPPFET W=1.16U L=0.12U M=1 
X15 net99 nmin2 net54 VDD LPPFET W=0.96U L=0.12U M=1 
X16 net87 B nmin1 VSS LPNFET W=0.86U L=0.12U M=1 
X17 net87 nmin2 net54 VSS LPNFET W=0.68U L=0.12U M=1 
X18 net93 C net99 VSS LPNFET W=0.74U L=0.12U M=1 
X19 net93 nmin3 net87 VSS LPNFET W=0.68U L=0.12U M=1 
X2 VDD net93 Y VDD LPPFET W=1.3U L=0.12U M=1 
X20 net99 nmin2 nmin1 VSS LPNFET W=0.92U L=0.12U M=1 
X21 net99 B net54 VSS LPNFET W=0.68U L=0.12U M=1 
X3 Y net93 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X4 VDD C nmin3 VDD LPPFET W=0.42U L=0.12U M=1 
X5 nmin3 C VSS VSS LPNFET W=0.3U L=0.12U M=1 
X6 VDD B nmin2 VDD LPPFET W=0.94U L=0.12U M=1 
X7 nmin2 B VSS VSS LPNFET W=0.68U L=0.12U M=1 
X8 VDD A nmin1 VDD LPPFET W=1.28U L=0.12U M=1 
X9 nmin1 A VSS VSS LPNFET W=0.92U L=0.12U M=1 
.ENDS XNOR3X2TS 

**** 
*.SUBCKT XNOR3X4TS Y A B C 
.SUBCKT XNOR3X4TS Y A B C VSS VDD
X0 VDD nmin1 net54 VDD LPPFET W=1.86U L=0.12U M=1 
X1 net54 nmin1 VSS VSS LPNFET W=1.48U L=0.12U M=1 
X10 net87 nmin2 nmin1 VDD LPPFET W=1.28U L=0.12U M=1 
X11 net87 B net54 VDD LPPFET W=2.06U L=0.12U M=1 
X12 net93 nmin3 net99 VDD LPPFET W=1.84U L=0.12U M=1 
X13 net93 C net87 VDD LPPFET W=1.84U L=0.12U M=1 
X14 net99 B nmin1 VDD LPPFET W=1.18U L=0.12U M=1 
X15 net99 nmin2 net54 VDD LPPFET W=1.8U L=0.12U M=1 
X16 net87 B nmin1 VSS LPNFET W=0.82U L=0.12U M=1 
X17 net87 nmin2 net54 VSS LPNFET W=1.42U L=0.12U M=1 
X18 net93 C net99 VSS LPNFET W=1.34U L=0.12U M=1 
X19 net93 nmin3 net87 VSS LPNFET W=1.38U L=0.12U M=1 
X2 VDD net93 Y VDD LPPFET W=2.6U L=0.12U M=1 
X20 net99 nmin2 nmin1 VSS LPNFET W=0.92U L=0.12U M=1 
X21 net99 B net54 VSS LPNFET W=1.42U L=0.12U M=1 
X3 Y net93 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X4 VDD C nmin3 VDD LPPFET W=0.84U L=0.12U M=1 
X5 nmin3 C VSS VSS LPNFET W=0.6U L=0.12U M=1 
X6 VDD B nmin2 VDD LPPFET W=1.12U L=0.12U M=1 
X7 nmin2 B VSS VSS LPNFET W=0.82U L=0.12U M=1 
X8 VDD A nmin1 VDD LPPFET W=1.28U L=0.12U M=1 
X9 nmin1 A VSS VSS LPNFET W=0.92U L=0.12U M=1 
.ENDS XNOR3X4TS 

**** 
*.SUBCKT XNOR3XLTS Y A B C 
.SUBCKT XNOR3XLTS Y A B C VSS VDD
X0 VDD nmin1 net54 VDD LPPFET W=0.28U L=0.12U M=1 
X1 net54 nmin1 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X10 net87 nmin2 nmin1 VDD LPPFET W=0.28U L=0.12U M=1 
X11 net87 B net54 VDD LPPFET W=0.28U L=0.12U M=1 
X12 net93 nmin3 net99 VDD LPPFET W=0.28U L=0.12U M=1 
X13 net93 C net87 VDD LPPFET W=0.28U L=0.12U M=1 
X14 net99 B nmin1 VDD LPPFET W=0.28U L=0.12U M=1 
X15 net99 nmin2 net54 VDD LPPFET W=0.28U L=0.12U M=1 
X16 net87 B nmin1 VSS LPNFET W=0.2U L=0.12U M=1 
X17 net87 nmin2 net54 VSS LPNFET W=0.2U L=0.12U M=1 
X18 net93 C net99 VSS LPNFET W=0.2U L=0.12U M=1 
X19 net93 nmin3 net87 VSS LPNFET W=0.2U L=0.12U M=1 
X2 VDD net93 Y VDD LPPFET W=0.42U L=0.12U M=1 
X20 net99 nmin2 nmin1 VSS LPNFET W=0.2U L=0.12U M=1 
X21 net99 B net54 VSS LPNFET W=0.2U L=0.12U M=1 
X3 Y net93 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X4 VDD C nmin3 VDD LPPFET W=0.28U L=0.12U M=1 
X5 nmin3 C VSS VSS LPNFET W=0.2U L=0.12U M=1 
X6 VDD B nmin2 VDD LPPFET W=0.28U L=0.12U M=1 
X7 nmin2 B VSS VSS LPNFET W=0.2U L=0.12U M=1 
X8 VDD A nmin1 VDD LPPFET W=0.28U L=0.12U M=1 
X9 nmin1 A VSS VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS XNOR3XLTS 

**** 
*.SUBCKT XOR2X1TS Y A B 
.SUBCKT XOR2X1TS Y A B VSS VDD
X0 Y A net35 VDD LPPFET W=0.76U L=0.12U M=1 
X1 Y nmin1 nmin2 VDD LPPFET W=0.78U L=0.12U M=1 
X2 Y nmin1 net35 VSS LPNFET W=0.56U L=0.12U M=1 
X3 Y A nmin2 VSS LPNFET W=0.54U L=0.12U M=1 
X4 VDD A nmin1 VDD LPPFET W=0.3U L=0.12U M=1 
X5 nmin1 A VSS VSS LPNFET W=0.22U L=0.12U M=1 
X6 VDD nmin2 net35 VDD LPPFET W=0.76U L=0.12U M=1 
X7 net35 nmin2 VSS VSS LPNFET W=0.56U L=0.12U M=1 
X8 VDD B nmin2 VDD LPPFET W=0.78U L=0.12U M=1 
X9 nmin2 B VSS VSS LPNFET W=0.54U L=0.12U M=1 
.ENDS XOR2X1TS 

**** 
*.SUBCKT XOR2X2TS Y A B 
.SUBCKT XOR2X2TS Y A B VSS VDD
X0 Y A net35 VDD LPPFET W=1.56U L=0.12U M=1 
X1 Y nmin1 nmin2 VDD LPPFET W=1.56U L=0.12U M=1 
X2 Y nmin1 net35 VSS LPNFET W=1.1U L=0.12U M=1 
X3 Y A nmin2 VSS LPNFET W=1.08U L=0.12U M=1 
X4 VDD A nmin1 VDD LPPFET W=0.62U L=0.12U M=1 
X5 nmin1 A VSS VSS LPNFET W=0.44U L=0.12U M=1 
X6 VDD nmin2 net35 VDD LPPFET W=1.56U L=0.12U M=1 
X7 net35 nmin2 VSS VSS LPNFET W=1.1U L=0.12U M=1 
X8 VDD B nmin2 VDD LPPFET W=1.56U L=0.12U M=1 
X9 nmin2 B VSS VSS LPNFET W=1.1U L=0.12U M=1 
.ENDS XOR2X2TS 

**** 
*.SUBCKT XOR2X4TS Y A B 
.SUBCKT XOR2X4TS Y A B VSS VDD
X0 Y A net35 VDD LPPFET W=3.12U L=0.12U M=1 
X1 Y nmin1 nmin2 VDD LPPFET W=3.12U L=0.12U M=1 
X2 Y nmin1 net35 VSS LPNFET W=2.16U L=0.12U M=1 
X3 Y A nmin2 VSS LPNFET W=2.16U L=0.12U M=1 
X4 VDD A nmin1 VDD LPPFET W=1.22U L=0.12U M=1 
X5 nmin1 A VSS VSS LPNFET W=0.88U L=0.12U M=1 
X6 VDD nmin2 net35 VDD LPPFET W=3.06U L=0.12U M=1 
X7 net35 nmin2 VSS VSS LPNFET W=2.16U L=0.12U M=1 
X8 VDD B nmin2 VDD LPPFET W=3.12U L=0.12U M=1 
X9 nmin2 B VSS VSS LPNFET W=2.2U L=0.12U M=1 
.ENDS XOR2X4TS 

**** 
*.SUBCKT XOR2XLTS Y A B 
.SUBCKT XOR2XLTS Y A B VSS VDD
X0 Y A net35 VDD LPPFET W=0.4U L=0.12U M=1 
X1 Y nmin1 nmin2 VDD LPPFET W=0.38U L=0.12U M=1 
X2 Y nmin1 net35 VSS LPNFET W=0.26U L=0.12U M=1 
X3 Y A nmin2 VSS LPNFET W=0.28U L=0.12U M=1 
X4 VDD A nmin1 VDD LPPFET W=0.28U L=0.12U M=1 
X5 nmin1 A VSS VSS LPNFET W=0.2U L=0.12U M=1 
X6 VDD nmin2 net35 VDD LPPFET W=0.4U L=0.12U M=1 
X7 net35 nmin2 VSS VSS LPNFET W=0.28U L=0.12U M=1 
X8 VDD B nmin2 VDD LPPFET W=0.4U L=0.12U M=1 
X9 nmin2 B VSS VSS LPNFET W=0.28U L=0.12U M=1 
.ENDS XOR2XLTS 

**** 
*.SUBCKT XOR3X1TS Y A B C 
.SUBCKT XOR3X1TS Y A B C VSS VDD
X0 VDD nmin1 net53 VDD LPPFET W=0.5U L=0.12U M=1 
X1 net53 nmin1 VSS VSS LPNFET W=0.36U L=0.12U M=1 
X10 net86 nmin2 nmin1 VDD LPPFET W=0.72U L=0.12U M=1 
X11 net86 B net53 VDD LPPFET W=0.5U L=0.12U M=1 
X12 net92 C net98 VDD LPPFET W=0.5U L=0.12U M=1 
X13 net92 nmin3 net86 VDD LPPFET W=0.5U L=0.12U M=1 
X14 net98 B nmin1 VDD LPPFET W=0.72U L=0.12U M=1 
X15 net98 nmin2 net53 VDD LPPFET W=0.5U L=0.12U M=1 
X16 net86 B nmin1 VSS LPNFET W=0.52U L=0.12U M=1 
X17 net86 nmin2 net53 VSS LPNFET W=0.36U L=0.12U M=1 
X18 net92 nmin3 net98 VSS LPNFET W=0.36U L=0.12U M=1 
X19 net92 C net86 VSS LPNFET W=0.36U L=0.12U M=1 
X2 VDD net92 Y VDD LPPFET W=0.64U L=0.12U M=1 
X20 net98 nmin2 nmin1 VSS LPNFET W=0.52U L=0.12U M=1 
X21 net98 B net53 VSS LPNFET W=0.36U L=0.12U M=1 
X3 Y net92 VSS VSS LPNFET W=0.46U L=0.12U M=1 
X4 VDD C nmin3 VDD LPPFET W=0.28U L=0.12U M=1 
X5 nmin3 C VSS VSS LPNFET W=0.2U L=0.12U M=1 
X6 VDD B nmin2 VDD LPPFET W=0.5U L=0.12U M=1 
X7 nmin2 B VSS VSS LPNFET W=0.36U L=0.12U M=1 
X8 VDD A nmin1 VDD LPPFET W=0.72U L=0.12U M=1 
X9 nmin1 A VSS VSS LPNFET W=0.52U L=0.12U M=1 
.ENDS XOR3X1TS 

**** 
*.SUBCKT XOR3X2TS Y A B C 
.SUBCKT XOR3X2TS Y A B C VSS VDD
X0 VDD nmin1 net53 VDD LPPFET W=0.96U L=0.12U M=1 
X1 net53 nmin1 VSS VSS LPNFET W=0.6U L=0.12U M=1 
X10 net86 nmin2 nmin1 VDD LPPFET W=1.28U L=0.12U M=1 
X11 net86 B net53 VDD LPPFET W=1.02U L=0.12U M=1 
X12 net92 C net98 VDD LPPFET W=0.98U L=0.12U M=1 
X13 net92 nmin3 net86 VDD LPPFET W=1.02U L=0.12U M=1 
X14 net98 B nmin1 VDD LPPFET W=1.16U L=0.12U M=1 
X15 net98 nmin2 net53 VDD LPPFET W=0.96U L=0.12U M=1 
X16 net86 B nmin1 VSS LPNFET W=0.86U L=0.12U M=1 
X17 net86 nmin2 net53 VSS LPNFET W=0.68U L=0.12U M=1 
X18 net92 nmin3 net98 VSS LPNFET W=0.68U L=0.12U M=1 
X19 net92 C net86 VSS LPNFET W=0.68U L=0.12U M=1 
X2 VDD net92 Y VDD LPPFET W=1.3U L=0.12U M=1 
X20 net98 nmin2 nmin1 VSS LPNFET W=0.92U L=0.12U M=1 
X21 net98 B net53 VSS LPNFET W=0.68U L=0.12U M=1 
X3 Y net92 VSS VSS LPNFET W=0.92U L=0.12U M=1 
X4 VDD C nmin3 VDD LPPFET W=0.42U L=0.12U M=1 
X5 nmin3 C VSS VSS LPNFET W=0.3U L=0.12U M=1 
X6 VDD B nmin2 VDD LPPFET W=0.94U L=0.12U M=1 
X7 nmin2 B VSS VSS LPNFET W=0.68U L=0.12U M=1 
X8 VDD A nmin1 VDD LPPFET W=1.28U L=0.12U M=1 
X9 nmin1 A VSS VSS LPNFET W=0.92U L=0.12U M=1 
.ENDS XOR3X2TS 

**** 
*.SUBCKT XOR3X4TS Y A B C 
.SUBCKT XOR3X4TS Y A B C VSS VDD
X0 VDD nmin1 net53 VDD LPPFET W=1.86U L=0.12U M=1 
X1 net53 nmin1 VSS VSS LPNFET W=1.48U L=0.12U M=1 
X10 net86 nmin2 nmin1 VDD LPPFET W=1.28U L=0.12U M=1 
X11 net86 B net53 VDD LPPFET W=2.06U L=0.12U M=1 
X12 net92 C net98 VDD LPPFET W=1.94U L=0.12U M=1 
X13 net92 nmin3 net86 VDD LPPFET W=2.06U L=0.12U M=1 
X14 net98 B nmin1 VDD LPPFET W=1.18U L=0.12U M=1 
X15 net98 nmin2 net53 VDD LPPFET W=1.8U L=0.12U M=1 
X16 net86 B nmin1 VSS LPNFET W=0.82U L=0.12U M=1 
X17 net86 nmin2 net53 VSS LPNFET W=1.42U L=0.12U M=1 
X18 net92 nmin3 net98 VSS LPNFET W=1.2U L=0.12U M=1 
X19 net92 C net86 VSS LPNFET W=1.48U L=0.12U M=1 
X2 VDD net92 Y VDD LPPFET W=2.6U L=0.12U M=1 
X20 net98 nmin2 nmin1 VSS LPNFET W=0.92U L=0.12U M=1 
X21 net98 B net53 VSS LPNFET W=1.42U L=0.12U M=1 
X3 Y net92 VSS VSS LPNFET W=1.84U L=0.12U M=1 
X4 VDD C nmin3 VDD LPPFET W=0.84U L=0.12U M=1 
X5 nmin3 C VSS VSS LPNFET W=0.6U L=0.12U M=1 
X6 VDD B nmin2 VDD LPPFET W=1.12U L=0.12U M=1 
X7 nmin2 B VSS VSS LPNFET W=0.82U L=0.12U M=1 
X8 VDD A nmin1 VDD LPPFET W=1.28U L=0.12U M=1 
X9 nmin1 A VSS VSS LPNFET W=0.92U L=0.12U M=1 
.ENDS XOR3X4TS 

**** 
*.SUBCKT XOR3XLTS Y A B C 
.SUBCKT XOR3XLTS Y A B C VSS VDD
X0 VDD nmin1 net53 VDD LPPFET W=0.28U L=0.12U M=1 
X1 net53 nmin1 VSS VSS LPNFET W=0.2U L=0.12U M=1 
X10 net86 nmin2 nmin1 VDD LPPFET W=0.28U L=0.12U M=1 
X11 net86 B net53 VDD LPPFET W=0.28U L=0.12U M=1 
X12 net92 C net98 VDD LPPFET W=0.28U L=0.12U M=1 
X13 net92 nmin3 net86 VDD LPPFET W=0.28U L=0.12U M=1 
X14 net98 B nmin1 VDD LPPFET W=0.28U L=0.12U M=1 
X15 net98 nmin2 net53 VDD LPPFET W=0.28U L=0.12U M=1 
X16 net86 B nmin1 VSS LPNFET W=0.2U L=0.12U M=1 
X17 net86 nmin2 net53 VSS LPNFET W=0.2U L=0.12U M=1 
X18 net92 nmin3 net98 VSS LPNFET W=0.2U L=0.12U M=1 
X19 net92 C net86 VSS LPNFET W=0.2U L=0.12U M=1 
X2 VDD net92 Y VDD LPPFET W=0.42U L=0.12U M=1 
X20 net98 nmin2 nmin1 VSS LPNFET W=0.2U L=0.12U M=1 
X21 net98 B net53 VSS LPNFET W=0.2U L=0.12U M=1 
X3 Y net92 VSS VSS LPNFET W=0.24U L=0.12U M=1 
X4 VDD C nmin3 VDD LPPFET W=0.28U L=0.12U M=1 
X5 nmin3 C VSS VSS LPNFET W=0.2U L=0.12U M=1 
X6 VDD B nmin2 VDD LPPFET W=0.28U L=0.12U M=1 
X7 nmin2 B VSS VSS LPNFET W=0.2U L=0.12U M=1 
X8 VDD A nmin1 VDD LPPFET W=0.28U L=0.12U M=1 
X9 nmin1 A VSS VSS LPNFET W=0.2U L=0.12U M=1 
.ENDS XOR3XLTS 
