
module aes_addroundkey ( clk, ld_r, text_in_r, w0, w1, w2, w3, sa00, sa01, 
        sa02, sa03, sa10, sa11, sa12, sa13, sa20, sa21, sa22, sa23, sa30, sa31, 
        sa32, sa33, sa00_next, sa01_next, sa02_next, sa03_next, sa10_next, 
        sa11_next, sa12_next, sa13_next, sa20_next, sa21_next, sa22_next, 
        sa23_next, sa30_next, sa31_next, sa32_next, sa33_next );
  input [127:0] text_in_r;
  input [31:0] w0;
  input [31:0] w1;
  input [31:0] w2;
  input [31:0] w3;
  output [7:0] sa00;
  output [7:0] sa01;
  output [7:0] sa02;
  output [7:0] sa03;
  output [7:0] sa10;
  output [7:0] sa11;
  output [7:0] sa12;
  output [7:0] sa13;
  output [7:0] sa20;
  output [7:0] sa21;
  output [7:0] sa22;
  output [7:0] sa23;
  output [7:0] sa30;
  output [7:0] sa31;
  output [7:0] sa32;
  output [7:0] sa33;
  input [7:0] sa00_next;
  input [7:0] sa01_next;
  input [7:0] sa02_next;
  input [7:0] sa03_next;
  input [7:0] sa10_next;
  input [7:0] sa11_next;
  input [7:0] sa12_next;
  input [7:0] sa13_next;
  input [7:0] sa20_next;
  input [7:0] sa21_next;
  input [7:0] sa22_next;
  input [7:0] sa23_next;
  input [7:0] sa30_next;
  input [7:0] sa31_next;
  input [7:0] sa32_next;
  input [7:0] sa33_next;
  input clk, ld_r;
  wire   \ux33/n10 , \ux33/n9 , \ux33/n8 , \ux33/n7 , \ux33/n6 , \ux33/n5 ,
         \ux33/n4 , \ux33/n3 , \ux33/n2 , \ux00/n18 , \ux00/n17 , \ux00/n16 ,
         \ux00/n15 , \ux00/n14 , \ux00/n13 , \ux00/n12 , \ux00/n11 ,
         \ux10/n18 , \ux10/n17 , \ux10/n16 , \ux10/n15 , \ux10/n14 ,
         \ux10/n13 , \ux10/n12 , \ux10/n11 , \ux20/n18 , \ux20/n17 ,
         \ux20/n16 , \ux20/n15 , \ux20/n14 , \ux20/n13 , \ux20/n12 ,
         \ux20/n11 , \ux30/n18 , \ux30/n17 , \ux30/n16 , \ux30/n15 ,
         \ux30/n14 , \ux30/n13 , \ux30/n12 , \ux30/n11 , \ux01/n18 ,
         \ux01/n17 , \ux01/n16 , \ux01/n15 , \ux01/n14 , \ux01/n13 ,
         \ux01/n12 , \ux01/n11 , \ux11/n18 , \ux11/n17 , \ux11/n16 ,
         \ux11/n15 , \ux11/n14 , \ux11/n13 , \ux11/n12 , \ux11/n11 ,
         \ux21/n18 , \ux21/n17 , \ux21/n16 , \ux21/n15 , \ux21/n14 ,
         \ux21/n13 , \ux21/n12 , \ux21/n11 , \ux31/n18 , \ux31/n17 ,
         \ux31/n16 , \ux31/n15 , \ux31/n14 , \ux31/n13 , \ux31/n12 ,
         \ux31/n11 , \ux02/n18 , \ux02/n17 , \ux02/n16 , \ux02/n15 ,
         \ux02/n14 , \ux02/n13 , \ux02/n12 , \ux02/n11 , \ux12/n18 ,
         \ux12/n17 , \ux12/n16 , \ux12/n15 , \ux12/n14 , \ux12/n13 ,
         \ux12/n12 , \ux12/n11 , \ux22/n18 , \ux22/n17 , \ux22/n16 ,
         \ux22/n15 , \ux22/n14 , \ux22/n13 , \ux22/n12 , \ux22/n11 ,
         \ux32/n18 , \ux32/n17 , \ux32/n16 , \ux32/n15 , \ux32/n14 ,
         \ux32/n13 , \ux32/n12 , \ux32/n11 , \ux03/n18 , \ux03/n17 ,
         \ux03/n16 , \ux03/n15 , \ux03/n14 , \ux03/n13 , \ux03/n12 ,
         \ux03/n11 , \ux13/n18 , \ux13/n17 , \ux13/n16 , \ux13/n15 ,
         \ux13/n14 , \ux13/n13 , \ux13/n12 , \ux13/n11 , \ux23/n18 ,
         \ux23/n17 , \ux23/n16 , \ux23/n15 , \ux23/n14 , \ux23/n13 ,
         \ux23/n12 , \ux23/n11 , n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080;
  assign \ux33/n10  = ld_r;

  SDFFQXLTS \ux33/sa_o_reg[0]  ( .D(sa33_next[0]), .SI(\ux33/n9 ), .SE(n1075), 
        .CK(clk), .Q(sa33[0]) );
  SDFFQXLTS \ux33/sa_o_reg[1]  ( .D(sa33_next[1]), .SI(\ux33/n8 ), .SE(n1039), 
        .CK(clk), .Q(sa33[1]) );
  SDFFQXLTS \ux33/sa_o_reg[2]  ( .D(sa33_next[2]), .SI(\ux33/n7 ), .SE(n1039), 
        .CK(clk), .Q(sa33[2]) );
  SDFFQXLTS \ux33/sa_o_reg[3]  ( .D(sa33_next[3]), .SI(\ux33/n6 ), .SE(n1039), 
        .CK(clk), .Q(sa33[3]) );
  SDFFQXLTS \ux33/sa_o_reg[4]  ( .D(sa33_next[4]), .SI(\ux33/n5 ), .SE(n1080), 
        .CK(clk), .Q(sa33[4]) );
  SDFFQXLTS \ux33/sa_o_reg[5]  ( .D(sa33_next[5]), .SI(\ux33/n4 ), .SE(n1069), 
        .CK(clk), .Q(sa33[5]) );
  SDFFQXLTS \ux33/sa_o_reg[6]  ( .D(sa33_next[6]), .SI(\ux33/n3 ), .SE(n1069), 
        .CK(clk), .Q(sa33[6]) );
  SDFFQXLTS \ux33/sa_o_reg[7]  ( .D(sa33_next[7]), .SI(\ux33/n2 ), .SE(n1080), 
        .CK(clk), .Q(sa33[7]) );
  SDFFQXLTS \ux00/sa_o_reg[0]  ( .D(sa00_next[0]), .SI(\ux00/n11 ), .SE(n1054), 
        .CK(clk), .Q(sa00[0]) );
  SDFFQXLTS \ux00/sa_o_reg[1]  ( .D(sa00_next[1]), .SI(\ux00/n12 ), .SE(n1053), 
        .CK(clk), .Q(sa00[1]) );
  SDFFQXLTS \ux00/sa_o_reg[2]  ( .D(sa00_next[2]), .SI(\ux00/n13 ), .SE(n1053), 
        .CK(clk), .Q(sa00[2]) );
  SDFFQXLTS \ux00/sa_o_reg[3]  ( .D(sa00_next[3]), .SI(\ux00/n14 ), .SE(n1053), 
        .CK(clk), .Q(sa00[3]) );
  SDFFQXLTS \ux00/sa_o_reg[4]  ( .D(sa00_next[4]), .SI(\ux00/n15 ), .SE(n1054), 
        .CK(clk), .Q(sa00[4]) );
  SDFFQXLTS \ux00/sa_o_reg[5]  ( .D(sa00_next[5]), .SI(\ux00/n16 ), .SE(n1054), 
        .CK(clk), .Q(sa00[5]) );
  SDFFQXLTS \ux00/sa_o_reg[6]  ( .D(sa00_next[6]), .SI(\ux00/n17 ), .SE(n1054), 
        .CK(clk), .Q(sa00[6]) );
  SDFFQXLTS \ux00/sa_o_reg[7]  ( .D(sa00_next[7]), .SI(\ux00/n18 ), .SE(n1055), 
        .CK(clk), .Q(sa00[7]) );
  SDFFQXLTS \ux10/sa_o_reg[0]  ( .D(sa10_next[0]), .SI(\ux10/n11 ), .SE(n1050), 
        .CK(clk), .Q(sa10[0]) );
  SDFFQXLTS \ux10/sa_o_reg[1]  ( .D(sa10_next[1]), .SI(\ux10/n12 ), .SE(n1049), 
        .CK(clk), .Q(sa10[1]) );
  SDFFQXLTS \ux10/sa_o_reg[2]  ( .D(sa10_next[2]), .SI(\ux10/n13 ), .SE(n1049), 
        .CK(clk), .Q(sa10[2]) );
  SDFFQXLTS \ux10/sa_o_reg[3]  ( .D(sa10_next[3]), .SI(\ux10/n14 ), .SE(n1049), 
        .CK(clk), .Q(sa10[3]) );
  SDFFQXLTS \ux10/sa_o_reg[4]  ( .D(sa10_next[4]), .SI(\ux10/n15 ), .SE(n1058), 
        .CK(clk), .Q(sa10[4]) );
  SDFFQXLTS \ux10/sa_o_reg[5]  ( .D(sa10_next[5]), .SI(\ux10/n16 ), .SE(n1058), 
        .CK(clk), .Q(sa10[5]) );
  SDFFQXLTS \ux10/sa_o_reg[6]  ( .D(sa10_next[6]), .SI(\ux10/n17 ), .SE(n1058), 
        .CK(clk), .Q(sa10[6]) );
  SDFFQXLTS \ux10/sa_o_reg[7]  ( .D(sa10_next[7]), .SI(\ux10/n18 ), .SE(n1059), 
        .CK(clk), .Q(sa10[7]) );
  SDFFQXLTS \ux20/sa_o_reg[0]  ( .D(sa20_next[0]), .SI(\ux20/n11 ), .SE(n1046), 
        .CK(clk), .Q(sa20[0]) );
  SDFFQXLTS \ux20/sa_o_reg[1]  ( .D(sa20_next[1]), .SI(\ux20/n12 ), .SE(n1045), 
        .CK(clk), .Q(sa20[1]) );
  SDFFQXLTS \ux20/sa_o_reg[2]  ( .D(sa20_next[2]), .SI(\ux20/n13 ), .SE(n1045), 
        .CK(clk), .Q(sa20[2]) );
  SDFFQXLTS \ux20/sa_o_reg[3]  ( .D(sa20_next[3]), .SI(\ux20/n14 ), .SE(n1045), 
        .CK(clk), .Q(sa20[3]) );
  SDFFQXLTS \ux20/sa_o_reg[4]  ( .D(sa20_next[4]), .SI(\ux20/n15 ), .SE(n1062), 
        .CK(clk), .Q(sa20[4]) );
  SDFFQXLTS \ux20/sa_o_reg[5]  ( .D(sa20_next[5]), .SI(\ux20/n16 ), .SE(n1062), 
        .CK(clk), .Q(sa20[5]) );
  SDFFQXLTS \ux20/sa_o_reg[6]  ( .D(sa20_next[6]), .SI(\ux20/n17 ), .SE(n1062), 
        .CK(clk), .Q(sa20[6]) );
  SDFFQXLTS \ux20/sa_o_reg[7]  ( .D(sa20_next[7]), .SI(\ux20/n18 ), .SE(n1063), 
        .CK(clk), .Q(sa20[7]) );
  SDFFQXLTS \ux30/sa_o_reg[0]  ( .D(sa30_next[0]), .SI(\ux30/n11 ), .SE(n1042), 
        .CK(clk), .Q(sa30[0]) );
  SDFFQXLTS \ux30/sa_o_reg[1]  ( .D(sa30_next[1]), .SI(\ux30/n12 ), .SE(n1041), 
        .CK(clk), .Q(sa30[1]) );
  SDFFQXLTS \ux30/sa_o_reg[2]  ( .D(sa30_next[2]), .SI(\ux30/n13 ), .SE(n1041), 
        .CK(clk), .Q(sa30[2]) );
  SDFFQXLTS \ux30/sa_o_reg[3]  ( .D(sa30_next[3]), .SI(\ux30/n14 ), .SE(n1041), 
        .CK(clk), .Q(sa30[3]) );
  SDFFQXLTS \ux30/sa_o_reg[4]  ( .D(sa30_next[4]), .SI(\ux30/n15 ), .SE(n1066), 
        .CK(clk), .Q(sa30[4]) );
  SDFFQXLTS \ux30/sa_o_reg[5]  ( .D(sa30_next[5]), .SI(\ux30/n16 ), .SE(n1066), 
        .CK(clk), .Q(sa30[5]) );
  SDFFQXLTS \ux30/sa_o_reg[6]  ( .D(sa30_next[6]), .SI(\ux30/n17 ), .SE(n1066), 
        .CK(clk), .Q(sa30[6]) );
  SDFFQXLTS \ux30/sa_o_reg[7]  ( .D(sa30_next[7]), .SI(\ux30/n18 ), .SE(n1066), 
        .CK(clk), .Q(sa30[7]) );
  SDFFQXLTS \ux01/sa_o_reg[0]  ( .D(sa01_next[0]), .SI(\ux01/n11 ), .SE(n1053), 
        .CK(clk), .Q(sa01[0]) );
  SDFFQXLTS \ux01/sa_o_reg[1]  ( .D(sa01_next[1]), .SI(\ux01/n12 ), .SE(n1052), 
        .CK(clk), .Q(sa01[1]) );
  SDFFQXLTS \ux01/sa_o_reg[2]  ( .D(sa01_next[2]), .SI(\ux01/n13 ), .SE(n1052), 
        .CK(clk), .Q(sa01[2]) );
  SDFFQXLTS \ux01/sa_o_reg[3]  ( .D(sa01_next[3]), .SI(\ux01/n14 ), .SE(n1052), 
        .CK(clk), .Q(sa01[3]) );
  SDFFQXLTS \ux01/sa_o_reg[4]  ( .D(sa01_next[4]), .SI(\ux01/n15 ), .SE(n1055), 
        .CK(clk), .Q(sa01[4]) );
  SDFFQXLTS \ux01/sa_o_reg[5]  ( .D(sa01_next[5]), .SI(\ux01/n16 ), .SE(n1055), 
        .CK(clk), .Q(sa01[5]) );
  SDFFQXLTS \ux01/sa_o_reg[6]  ( .D(sa01_next[6]), .SI(\ux01/n17 ), .SE(n1055), 
        .CK(clk), .Q(sa01[6]) );
  SDFFQXLTS \ux01/sa_o_reg[7]  ( .D(sa01_next[7]), .SI(\ux01/n18 ), .SE(n1056), 
        .CK(clk), .Q(sa01[7]) );
  SDFFQXLTS \ux11/sa_o_reg[0]  ( .D(sa11_next[0]), .SI(\ux11/n11 ), .SE(n1049), 
        .CK(clk), .Q(sa11[0]) );
  SDFFQXLTS \ux11/sa_o_reg[1]  ( .D(sa11_next[1]), .SI(\ux11/n12 ), .SE(n1048), 
        .CK(clk), .Q(sa11[1]) );
  SDFFQXLTS \ux11/sa_o_reg[2]  ( .D(sa11_next[2]), .SI(\ux11/n13 ), .SE(n1048), 
        .CK(clk), .Q(sa11[2]) );
  SDFFQXLTS \ux11/sa_o_reg[3]  ( .D(sa11_next[3]), .SI(\ux11/n14 ), .SE(n1048), 
        .CK(clk), .Q(sa11[3]) );
  SDFFQXLTS \ux11/sa_o_reg[4]  ( .D(sa11_next[4]), .SI(\ux11/n15 ), .SE(n1059), 
        .CK(clk), .Q(sa11[4]) );
  SDFFQXLTS \ux11/sa_o_reg[5]  ( .D(sa11_next[5]), .SI(\ux11/n16 ), .SE(n1059), 
        .CK(clk), .Q(sa11[5]) );
  SDFFQXLTS \ux11/sa_o_reg[6]  ( .D(sa11_next[6]), .SI(\ux11/n17 ), .SE(n1059), 
        .CK(clk), .Q(sa11[6]) );
  SDFFQXLTS \ux11/sa_o_reg[7]  ( .D(sa11_next[7]), .SI(\ux11/n18 ), .SE(n1060), 
        .CK(clk), .Q(sa11[7]) );
  SDFFQXLTS \ux21/sa_o_reg[0]  ( .D(sa21_next[0]), .SI(\ux21/n11 ), .SE(n1045), 
        .CK(clk), .Q(sa21[0]) );
  SDFFQXLTS \ux21/sa_o_reg[1]  ( .D(sa21_next[1]), .SI(\ux21/n12 ), .SE(n1044), 
        .CK(clk), .Q(sa21[1]) );
  SDFFQXLTS \ux21/sa_o_reg[2]  ( .D(sa21_next[2]), .SI(\ux21/n13 ), .SE(n1044), 
        .CK(clk), .Q(sa21[2]) );
  SDFFQXLTS \ux21/sa_o_reg[3]  ( .D(sa21_next[3]), .SI(\ux21/n14 ), .SE(n1044), 
        .CK(clk), .Q(sa21[3]) );
  SDFFQXLTS \ux21/sa_o_reg[4]  ( .D(sa21_next[4]), .SI(\ux21/n15 ), .SE(n1063), 
        .CK(clk), .Q(sa21[4]) );
  SDFFQXLTS \ux21/sa_o_reg[5]  ( .D(sa21_next[5]), .SI(\ux21/n16 ), .SE(n1063), 
        .CK(clk), .Q(sa21[5]) );
  SDFFQXLTS \ux21/sa_o_reg[6]  ( .D(sa21_next[6]), .SI(\ux21/n17 ), .SE(n1063), 
        .CK(clk), .Q(sa21[6]) );
  SDFFQXLTS \ux21/sa_o_reg[7]  ( .D(sa21_next[7]), .SI(\ux21/n18 ), .SE(n1064), 
        .CK(clk), .Q(sa21[7]) );
  SDFFQXLTS \ux31/sa_o_reg[0]  ( .D(sa31_next[0]), .SI(\ux31/n11 ), .SE(n1041), 
        .CK(clk), .Q(sa31[0]) );
  SDFFQXLTS \ux31/sa_o_reg[1]  ( .D(sa31_next[1]), .SI(\ux31/n12 ), .SE(n1040), 
        .CK(clk), .Q(sa31[1]) );
  SDFFQXLTS \ux31/sa_o_reg[2]  ( .D(sa31_next[2]), .SI(\ux31/n13 ), .SE(n1040), 
        .CK(clk), .Q(sa31[2]) );
  SDFFQXLTS \ux31/sa_o_reg[3]  ( .D(sa31_next[3]), .SI(\ux31/n14 ), .SE(n1040), 
        .CK(clk), .Q(sa31[3]) );
  SDFFQXLTS \ux31/sa_o_reg[4]  ( .D(sa31_next[4]), .SI(\ux31/n15 ), .SE(n1067), 
        .CK(clk), .Q(sa31[4]) );
  SDFFQXLTS \ux31/sa_o_reg[5]  ( .D(sa31_next[5]), .SI(\ux31/n16 ), .SE(n1067), 
        .CK(clk), .Q(sa31[5]) );
  SDFFQXLTS \ux31/sa_o_reg[6]  ( .D(sa31_next[6]), .SI(\ux31/n17 ), .SE(n1067), 
        .CK(clk), .Q(sa31[6]) );
  SDFFQXLTS \ux31/sa_o_reg[7]  ( .D(sa31_next[7]), .SI(\ux31/n18 ), .SE(n1067), 
        .CK(clk), .Q(sa31[7]) );
  SDFFQXLTS \ux02/sa_o_reg[0]  ( .D(sa02_next[0]), .SI(\ux02/n11 ), .SE(n1052), 
        .CK(clk), .Q(sa02[0]) );
  SDFFQXLTS \ux02/sa_o_reg[1]  ( .D(sa02_next[1]), .SI(\ux02/n12 ), .SE(n1051), 
        .CK(clk), .Q(sa02[1]) );
  SDFFQXLTS \ux02/sa_o_reg[2]  ( .D(sa02_next[2]), .SI(\ux02/n13 ), .SE(n1051), 
        .CK(clk), .Q(sa02[2]) );
  SDFFQXLTS \ux02/sa_o_reg[3]  ( .D(sa02_next[3]), .SI(\ux02/n14 ), .SE(n1051), 
        .CK(clk), .Q(sa02[3]) );
  SDFFQXLTS \ux02/sa_o_reg[4]  ( .D(sa02_next[4]), .SI(\ux02/n15 ), .SE(n1056), 
        .CK(clk), .Q(sa02[4]) );
  SDFFQXLTS \ux02/sa_o_reg[5]  ( .D(sa02_next[5]), .SI(\ux02/n16 ), .SE(n1056), 
        .CK(clk), .Q(sa02[5]) );
  SDFFQXLTS \ux02/sa_o_reg[6]  ( .D(sa02_next[6]), .SI(\ux02/n17 ), .SE(n1056), 
        .CK(clk), .Q(sa02[6]) );
  SDFFQXLTS \ux02/sa_o_reg[7]  ( .D(sa02_next[7]), .SI(\ux02/n18 ), .SE(n1057), 
        .CK(clk), .Q(sa02[7]) );
  SDFFQXLTS \ux12/sa_o_reg[0]  ( .D(sa12_next[0]), .SI(\ux12/n11 ), .SE(n1048), 
        .CK(clk), .Q(sa12[0]) );
  SDFFQXLTS \ux12/sa_o_reg[1]  ( .D(sa12_next[1]), .SI(\ux12/n12 ), .SE(n1047), 
        .CK(clk), .Q(sa12[1]) );
  SDFFQXLTS \ux12/sa_o_reg[2]  ( .D(sa12_next[2]), .SI(\ux12/n13 ), .SE(n1047), 
        .CK(clk), .Q(sa12[2]) );
  SDFFQXLTS \ux12/sa_o_reg[3]  ( .D(sa12_next[3]), .SI(\ux12/n14 ), .SE(n1047), 
        .CK(clk), .Q(sa12[3]) );
  SDFFQXLTS \ux12/sa_o_reg[4]  ( .D(sa12_next[4]), .SI(\ux12/n15 ), .SE(n1060), 
        .CK(clk), .Q(sa12[4]) );
  SDFFQXLTS \ux12/sa_o_reg[5]  ( .D(sa12_next[5]), .SI(\ux12/n16 ), .SE(n1060), 
        .CK(clk), .Q(sa12[5]) );
  SDFFQXLTS \ux12/sa_o_reg[6]  ( .D(sa12_next[6]), .SI(\ux12/n17 ), .SE(n1060), 
        .CK(clk), .Q(sa12[6]) );
  SDFFQXLTS \ux12/sa_o_reg[7]  ( .D(sa12_next[7]), .SI(\ux12/n18 ), .SE(n1061), 
        .CK(clk), .Q(sa12[7]) );
  SDFFQXLTS \ux22/sa_o_reg[0]  ( .D(sa22_next[0]), .SI(\ux22/n11 ), .SE(n1044), 
        .CK(clk), .Q(sa22[0]) );
  SDFFQXLTS \ux22/sa_o_reg[1]  ( .D(sa22_next[1]), .SI(\ux22/n12 ), .SE(n1043), 
        .CK(clk), .Q(sa22[1]) );
  SDFFQXLTS \ux22/sa_o_reg[2]  ( .D(sa22_next[2]), .SI(\ux22/n13 ), .SE(n1043), 
        .CK(clk), .Q(sa22[2]) );
  SDFFQXLTS \ux22/sa_o_reg[3]  ( .D(sa22_next[3]), .SI(\ux22/n14 ), .SE(n1043), 
        .CK(clk), .Q(sa22[3]) );
  SDFFQXLTS \ux22/sa_o_reg[4]  ( .D(sa22_next[4]), .SI(\ux22/n15 ), .SE(n1064), 
        .CK(clk), .Q(sa22[4]) );
  SDFFQXLTS \ux22/sa_o_reg[5]  ( .D(sa22_next[5]), .SI(\ux22/n16 ), .SE(n1064), 
        .CK(clk), .Q(sa22[5]) );
  SDFFQXLTS \ux22/sa_o_reg[6]  ( .D(sa22_next[6]), .SI(\ux22/n17 ), .SE(n1064), 
        .CK(clk), .Q(sa22[6]) );
  SDFFQXLTS \ux22/sa_o_reg[7]  ( .D(sa22_next[7]), .SI(\ux22/n18 ), .SE(n1065), 
        .CK(clk), .Q(sa22[7]) );
  SDFFQXLTS \ux32/sa_o_reg[0]  ( .D(sa32_next[0]), .SI(\ux32/n11 ), .SE(n1040), 
        .CK(clk), .Q(sa32[0]) );
  SDFFQXLTS \ux32/sa_o_reg[1]  ( .D(sa32_next[1]), .SI(\ux32/n12 ), .SE(n1073), 
        .CK(clk), .Q(sa32[1]) );
  SDFFQXLTS \ux32/sa_o_reg[2]  ( .D(sa32_next[2]), .SI(\ux32/n13 ), .SE(n1074), 
        .CK(clk), .Q(sa32[2]) );
  SDFFQXLTS \ux32/sa_o_reg[3]  ( .D(sa32_next[3]), .SI(\ux32/n14 ), .SE(n1078), 
        .CK(clk), .Q(sa32[3]) );
  SDFFQXLTS \ux32/sa_o_reg[4]  ( .D(sa32_next[4]), .SI(\ux32/n15 ), .SE(n1068), 
        .CK(clk), .Q(sa32[4]) );
  SDFFQXLTS \ux32/sa_o_reg[5]  ( .D(sa32_next[5]), .SI(\ux32/n16 ), .SE(n1068), 
        .CK(clk), .Q(sa32[5]) );
  SDFFQXLTS \ux32/sa_o_reg[6]  ( .D(sa32_next[6]), .SI(\ux32/n17 ), .SE(n1068), 
        .CK(clk), .Q(sa32[6]) );
  SDFFQXLTS \ux32/sa_o_reg[7]  ( .D(sa32_next[7]), .SI(\ux32/n18 ), .SE(n1068), 
        .CK(clk), .Q(sa32[7]) );
  SDFFQXLTS \ux03/sa_o_reg[0]  ( .D(sa03_next[0]), .SI(\ux03/n11 ), .SE(n1051), 
        .CK(clk), .Q(sa03[0]) );
  SDFFQXLTS \ux03/sa_o_reg[1]  ( .D(sa03_next[1]), .SI(\ux03/n12 ), .SE(n1050), 
        .CK(clk), .Q(sa03[1]) );
  SDFFQXLTS \ux03/sa_o_reg[2]  ( .D(sa03_next[2]), .SI(\ux03/n13 ), .SE(n1050), 
        .CK(clk), .Q(sa03[2]) );
  SDFFQXLTS \ux03/sa_o_reg[3]  ( .D(sa03_next[3]), .SI(\ux03/n14 ), .SE(n1050), 
        .CK(clk), .Q(sa03[3]) );
  SDFFQXLTS \ux03/sa_o_reg[4]  ( .D(sa03_next[4]), .SI(\ux03/n15 ), .SE(n1057), 
        .CK(clk), .Q(sa03[4]) );
  SDFFQXLTS \ux03/sa_o_reg[5]  ( .D(sa03_next[5]), .SI(\ux03/n16 ), .SE(n1057), 
        .CK(clk), .Q(sa03[5]) );
  SDFFQXLTS \ux03/sa_o_reg[6]  ( .D(sa03_next[6]), .SI(\ux03/n17 ), .SE(n1057), 
        .CK(clk), .Q(sa03[6]) );
  SDFFQXLTS \ux03/sa_o_reg[7]  ( .D(sa03_next[7]), .SI(\ux03/n18 ), .SE(n1058), 
        .CK(clk), .Q(sa03[7]) );
  SDFFQXLTS \ux13/sa_o_reg[0]  ( .D(sa13_next[0]), .SI(\ux13/n11 ), .SE(n1047), 
        .CK(clk), .Q(sa13[0]) );
  SDFFQXLTS \ux13/sa_o_reg[1]  ( .D(sa13_next[1]), .SI(\ux13/n12 ), .SE(n1046), 
        .CK(clk), .Q(sa13[1]) );
  SDFFQXLTS \ux13/sa_o_reg[2]  ( .D(sa13_next[2]), .SI(\ux13/n13 ), .SE(n1046), 
        .CK(clk), .Q(sa13[2]) );
  SDFFQXLTS \ux13/sa_o_reg[3]  ( .D(sa13_next[3]), .SI(\ux13/n14 ), .SE(n1046), 
        .CK(clk), .Q(sa13[3]) );
  SDFFQXLTS \ux13/sa_o_reg[4]  ( .D(sa13_next[4]), .SI(\ux13/n15 ), .SE(n1061), 
        .CK(clk), .Q(sa13[4]) );
  SDFFQXLTS \ux13/sa_o_reg[5]  ( .D(sa13_next[5]), .SI(\ux13/n16 ), .SE(n1061), 
        .CK(clk), .Q(sa13[5]) );
  SDFFQXLTS \ux13/sa_o_reg[6]  ( .D(sa13_next[6]), .SI(\ux13/n17 ), .SE(n1061), 
        .CK(clk), .Q(sa13[6]) );
  SDFFQXLTS \ux13/sa_o_reg[7]  ( .D(sa13_next[7]), .SI(\ux13/n18 ), .SE(n1062), 
        .CK(clk), .Q(sa13[7]) );
  SDFFQXLTS \ux23/sa_o_reg[0]  ( .D(sa23_next[0]), .SI(\ux23/n11 ), .SE(n1043), 
        .CK(clk), .Q(sa23[0]) );
  SDFFQXLTS \ux23/sa_o_reg[1]  ( .D(sa23_next[1]), .SI(\ux23/n12 ), .SE(n1042), 
        .CK(clk), .Q(sa23[1]) );
  SDFFQXLTS \ux23/sa_o_reg[2]  ( .D(sa23_next[2]), .SI(\ux23/n13 ), .SE(n1042), 
        .CK(clk), .Q(sa23[2]) );
  SDFFQXLTS \ux23/sa_o_reg[3]  ( .D(sa23_next[3]), .SI(\ux23/n14 ), .SE(n1042), 
        .CK(clk), .Q(sa23[3]) );
  SDFFQXLTS \ux23/sa_o_reg[4]  ( .D(sa23_next[4]), .SI(\ux23/n15 ), .SE(n1065), 
        .CK(clk), .Q(sa23[4]) );
  SDFFQXLTS \ux23/sa_o_reg[5]  ( .D(sa23_next[5]), .SI(\ux23/n16 ), .SE(n1065), 
        .CK(clk), .Q(sa23[5]) );
  SDFFQXLTS \ux23/sa_o_reg[6]  ( .D(sa23_next[6]), .SI(\ux23/n17 ), .SE(n1065), 
        .CK(clk), .Q(sa23[6]) );
  SDFFQXLTS \ux23/sa_o_reg[7]  ( .D(sa23_next[7]), .SI(\ux23/n18 ), .SE(n1039), 
        .CK(clk), .Q(sa23[7]) );
  XOR2X1TS U14 ( .A(n902), .B(n646), .Y(\ux32/n13 ) );
  XOR2X1TS U16 ( .A(n910), .B(n654), .Y(\ux32/n11 ) );
  XOR2X1TS U70 ( .A(n966), .B(n710), .Y(\ux13/n13 ) );
  XOR2X1TS U10 ( .A(n886), .B(n630), .Y(\ux32/n17 ) );
  XOR2X1TS U11 ( .A(n890), .B(n634), .Y(\ux32/n16 ) );
  XOR2X1TS U69 ( .A(n962), .B(n706), .Y(\ux13/n14 ) );
  XOR2X1TS U9 ( .A(n882), .B(n626), .Y(\ux32/n18 ) );
  XOR2X1TS U102 ( .A(n934), .B(n678), .Y(\ux03/n13 ) );
  XOR2X1TS U66 ( .A(n950), .B(n694), .Y(\ux13/n17 ) );
  XOR2X1TS U100 ( .A(n926), .B(n670), .Y(\ux03/n15 ) );
  XOR2X1TS U43 ( .A(n858), .B(n602), .Y(\ux22/n16 ) );
  XOR2X1TS U103 ( .A(n938), .B(n682), .Y(\ux03/n12 ) );
  XOR2X1TS U15 ( .A(n906), .B(n650), .Y(\ux32/n12 ) );
  XOR2X1TS U72 ( .A(n974), .B(n718), .Y(\ux13/n11 ) );
  XOR2X1TS U44 ( .A(n862), .B(n606), .Y(\ux22/n15 ) );
  XOR2X1TS U98 ( .A(n918), .B(n662), .Y(\ux03/n17 ) );
  XOR2X1TS U39 ( .A(n1002), .B(n746), .Y(\ux23/n12 ) );
  XOR2X1TS U71 ( .A(n970), .B(n714), .Y(\ux13/n12 ) );
  XOR2X1TS U45 ( .A(n866), .B(n610), .Y(\ux22/n14 ) );
  XOR2X1TS U99 ( .A(n922), .B(n666), .Y(\ux03/n16 ) );
  XOR2X1TS U41 ( .A(n850), .B(n594), .Y(\ux22/n18 ) );
  XOR2X1TS U37 ( .A(n994), .B(n738), .Y(\ux23/n14 ) );
  XOR2X1TS U46 ( .A(n870), .B(n614), .Y(\ux22/n13 ) );
  XOR2X1TS U97 ( .A(n914), .B(n658), .Y(\ux03/n18 ) );
  XOR2X1TS U42 ( .A(n854), .B(n598), .Y(\ux22/n17 ) );
  XOR2X1TS U104 ( .A(n942), .B(n686), .Y(\ux03/n11 ) );
  XOR2X1TS U47 ( .A(n874), .B(n618), .Y(\ux22/n12 ) );
  XOR2X1TS U13 ( .A(n898), .B(n642), .Y(\ux32/n14 ) );
  XOR2X1TS U36 ( .A(n990), .B(n734), .Y(\ux23/n15 ) );
  XOR2X1TS U65 ( .A(n946), .B(n690), .Y(\ux13/n18 ) );
  XOR2X1TS U48 ( .A(n878), .B(n622), .Y(\ux22/n11 ) );
  XOR2X1TS U35 ( .A(n986), .B(n730), .Y(\ux23/n16 ) );
  XOR2X1TS U68 ( .A(n958), .B(n702), .Y(\ux13/n15 ) );
  XOR2X1TS U40 ( .A(n1006), .B(n750), .Y(\ux23/n11 ) );
  XOR2X1TS U73 ( .A(n818), .B(n562), .Y(\ux12/n18 ) );
  XOR2X1TS U34 ( .A(n982), .B(n726), .Y(\ux23/n17 ) );
  XOR2X1TS U101 ( .A(n930), .B(n674), .Y(\ux03/n14 ) );
  XOR2X1TS U38 ( .A(n998), .B(n742), .Y(\ux23/n13 ) );
  XOR2X1TS U74 ( .A(n822), .B(n566), .Y(\ux12/n17 ) );
  XOR2X1TS U33 ( .A(n978), .B(n722), .Y(\ux23/n18 ) );
  XOR2X1TS U67 ( .A(n954), .B(n698), .Y(\ux13/n16 ) );
  XOR2X1TS U12 ( .A(n894), .B(n638), .Y(\ux32/n15 ) );
  XOR2X1TS U24 ( .A(n784), .B(n528), .Y(\ux31/n11 ) );
  XOR2X1TS U75 ( .A(n826), .B(n570), .Y(\ux12/n16 ) );
  XOR2X1TS U76 ( .A(n830), .B(n574), .Y(\ux12/n15 ) );
  XOR2X1TS U77 ( .A(n834), .B(n578), .Y(\ux12/n14 ) );
  XOR2X1TS U78 ( .A(n838), .B(n582), .Y(\ux12/n13 ) );
  XOR2X1TS U79 ( .A(n842), .B(n586), .Y(\ux12/n12 ) );
  XOR2X1TS U80 ( .A(n846), .B(n590), .Y(\ux12/n11 ) );
  XOR2X1TS U105 ( .A(n786), .B(n530), .Y(\ux02/n18 ) );
  XOR2X1TS U106 ( .A(n790), .B(n534), .Y(\ux02/n17 ) );
  XOR2X1TS U107 ( .A(n794), .B(n538), .Y(\ux02/n16 ) );
  XOR2X1TS U108 ( .A(n798), .B(n542), .Y(\ux02/n15 ) );
  XOR2X1TS U109 ( .A(n802), .B(n546), .Y(\ux02/n14 ) );
  XOR2X1TS U110 ( .A(n806), .B(n550), .Y(\ux02/n13 ) );
  XOR2X1TS U111 ( .A(n810), .B(n554), .Y(\ux02/n12 ) );
  XOR2X1TS U112 ( .A(n814), .B(n558), .Y(\ux02/n11 ) );
  XOR2X1TS U17 ( .A(n812), .B(n556), .Y(\ux31/n18 ) );
  XOR2X1TS U18 ( .A(n808), .B(n552), .Y(\ux31/n17 ) );
  XOR2X1TS U19 ( .A(n804), .B(n548), .Y(\ux31/n16 ) );
  XOR2X1TS U20 ( .A(n800), .B(n544), .Y(\ux31/n15 ) );
  XOR2X1TS U21 ( .A(n796), .B(n540), .Y(\ux31/n14 ) );
  XOR2X1TS U22 ( .A(n792), .B(n536), .Y(\ux31/n13 ) );
  XOR2X1TS U23 ( .A(n788), .B(n532), .Y(\ux31/n12 ) );
  XOR2X1TS U1 ( .A(n1038), .B(n782), .Y(\ux33/n9 ) );
  XOR2X1TS U49 ( .A(n844), .B(n588), .Y(\ux21/n18 ) );
  XOR2X1TS U50 ( .A(n840), .B(n584), .Y(\ux21/n17 ) );
  XOR2X1TS U51 ( .A(n836), .B(n580), .Y(\ux21/n16 ) );
  XOR2X1TS U52 ( .A(n832), .B(n576), .Y(\ux21/n15 ) );
  XOR2X1TS U53 ( .A(n828), .B(n572), .Y(\ux21/n14 ) );
  XOR2X1TS U54 ( .A(n824), .B(n568), .Y(\ux21/n13 ) );
  XOR2X1TS U55 ( .A(n820), .B(n564), .Y(\ux21/n12 ) );
  XOR2X1TS U56 ( .A(n816), .B(n560), .Y(\ux21/n11 ) );
  XOR2X1TS U81 ( .A(n876), .B(n620), .Y(\ux11/n18 ) );
  XOR2X1TS U82 ( .A(n872), .B(n616), .Y(\ux11/n17 ) );
  XOR2X1TS U83 ( .A(n868), .B(n612), .Y(\ux11/n16 ) );
  XOR2X1TS U84 ( .A(n864), .B(n608), .Y(\ux11/n15 ) );
  XOR2X1TS U85 ( .A(n860), .B(n604), .Y(\ux11/n14 ) );
  XOR2X1TS U86 ( .A(n856), .B(n600), .Y(\ux11/n13 ) );
  XOR2X1TS U87 ( .A(n852), .B(n596), .Y(\ux11/n12 ) );
  XOR2X1TS U88 ( .A(n848), .B(n592), .Y(\ux11/n11 ) );
  XOR2X1TS U113 ( .A(n908), .B(n652), .Y(\ux01/n18 ) );
  XOR2X1TS U114 ( .A(n904), .B(n648), .Y(\ux01/n17 ) );
  XOR2X1TS U115 ( .A(n900), .B(n644), .Y(\ux01/n16 ) );
  XOR2X1TS U116 ( .A(n896), .B(n640), .Y(\ux01/n15 ) );
  XOR2X1TS U117 ( .A(n892), .B(n636), .Y(\ux01/n14 ) );
  XOR2X1TS U118 ( .A(n888), .B(n632), .Y(\ux01/n13 ) );
  XOR2X1TS U119 ( .A(n884), .B(n628), .Y(\ux01/n12 ) );
  XOR2X1TS U120 ( .A(n880), .B(n624), .Y(\ux01/n11 ) );
  XOR2X1TS U25 ( .A(n940), .B(n684), .Y(\ux30/n18 ) );
  XOR2X1TS U26 ( .A(n936), .B(n680), .Y(\ux30/n17 ) );
  XOR2X1TS U27 ( .A(n932), .B(n676), .Y(\ux30/n16 ) );
  XOR2X1TS U28 ( .A(n928), .B(n672), .Y(\ux30/n15 ) );
  XOR2X1TS U29 ( .A(n924), .B(n668), .Y(\ux30/n14 ) );
  XOR2X1TS U30 ( .A(n920), .B(n664), .Y(\ux30/n13 ) );
  XOR2X1TS U31 ( .A(n916), .B(n660), .Y(\ux30/n12 ) );
  XOR2X1TS U32 ( .A(n912), .B(n656), .Y(\ux30/n11 ) );
  XOR2X1TS U57 ( .A(n972), .B(n716), .Y(\ux20/n18 ) );
  XOR2X1TS U58 ( .A(n968), .B(n712), .Y(\ux20/n17 ) );
  XOR2X1TS U59 ( .A(n964), .B(n708), .Y(\ux20/n16 ) );
  XOR2X1TS U60 ( .A(n960), .B(n704), .Y(\ux20/n15 ) );
  XOR2X1TS U61 ( .A(n956), .B(n700), .Y(\ux20/n14 ) );
  XOR2X1TS U62 ( .A(n952), .B(n696), .Y(\ux20/n13 ) );
  XOR2X1TS U63 ( .A(n948), .B(n692), .Y(\ux20/n12 ) );
  XOR2X1TS U64 ( .A(n944), .B(n688), .Y(\ux20/n11 ) );
  XOR2X1TS U89 ( .A(n1004), .B(n748), .Y(\ux10/n18 ) );
  XOR2X1TS U90 ( .A(n1000), .B(n744), .Y(\ux10/n17 ) );
  XOR2X1TS U91 ( .A(n996), .B(n740), .Y(\ux10/n16 ) );
  XOR2X1TS U92 ( .A(n992), .B(n736), .Y(\ux10/n15 ) );
  XOR2X1TS U93 ( .A(n988), .B(n732), .Y(\ux10/n14 ) );
  XOR2X1TS U94 ( .A(n984), .B(n728), .Y(\ux10/n13 ) );
  XOR2X1TS U95 ( .A(n980), .B(n724), .Y(\ux10/n12 ) );
  XOR2X1TS U96 ( .A(n976), .B(n720), .Y(\ux10/n11 ) );
  XOR2X1TS U121 ( .A(n1036), .B(n780), .Y(\ux00/n18 ) );
  XOR2X1TS U122 ( .A(n1032), .B(n776), .Y(\ux00/n17 ) );
  XOR2X1TS U123 ( .A(n1028), .B(n772), .Y(\ux00/n16 ) );
  XOR2X1TS U124 ( .A(n1024), .B(n768), .Y(\ux00/n15 ) );
  XOR2X1TS U125 ( .A(n1020), .B(n764), .Y(\ux00/n14 ) );
  XOR2X1TS U126 ( .A(n1016), .B(n760), .Y(\ux00/n13 ) );
  XOR2X1TS U127 ( .A(n1012), .B(n756), .Y(\ux00/n12 ) );
  XOR2X1TS U128 ( .A(n1008), .B(n752), .Y(\ux00/n11 ) );
  XOR2X1TS U8 ( .A(n1010), .B(n754), .Y(\ux33/n2 ) );
  XOR2X1TS U7 ( .A(n1014), .B(n758), .Y(\ux33/n3 ) );
  XOR2X1TS U6 ( .A(n1018), .B(n762), .Y(\ux33/n4 ) );
  XOR2X1TS U5 ( .A(n1022), .B(n766), .Y(\ux33/n5 ) );
  XOR2X1TS U4 ( .A(n1026), .B(n770), .Y(\ux33/n6 ) );
  XOR2X1TS U3 ( .A(n1030), .B(n774), .Y(\ux33/n7 ) );
  XOR2X1TS U2 ( .A(n1034), .B(n778), .Y(\ux33/n8 ) );
  CLKBUFX2TS U129 ( .A(n1079), .Y(n1071) );
  CLKBUFX2TS U130 ( .A(n1079), .Y(n1072) );
  CLKBUFX2TS U131 ( .A(n1069), .Y(n1068) );
  CLKBUFX2TS U132 ( .A(n1077), .Y(n1078) );
  CLKBUFX2TS U133 ( .A(n1078), .Y(n1074) );
  CLKBUFX2TS U134 ( .A(n1078), .Y(n1073) );
  CLKBUFX2TS U135 ( .A(n1070), .Y(n1065) );
  CLKBUFX2TS U136 ( .A(n1070), .Y(n1043) );
  CLKBUFX2TS U137 ( .A(n1071), .Y(n1061) );
  CLKBUFX2TS U138 ( .A(n1075), .Y(n1047) );
  CLKBUFX2TS U139 ( .A(n1072), .Y(n1057) );
  CLKBUFX2TS U140 ( .A(n1074), .Y(n1051) );
  CLKBUFX2TS U141 ( .A(n1069), .Y(n1067) );
  CLKBUFX2TS U142 ( .A(n1070), .Y(n1064) );
  CLKBUFX2TS U143 ( .A(n1071), .Y(n1044) );
  CLKBUFX2TS U144 ( .A(n1072), .Y(n1060) );
  CLKBUFX2TS U145 ( .A(n1075), .Y(n1048) );
  CLKBUFX2TS U146 ( .A(n1079), .Y(n1056) );
  CLKBUFX2TS U147 ( .A(n1073), .Y(n1052) );
  CLKBUFX2TS U148 ( .A(n1070), .Y(n1066) );
  CLKBUFX2TS U149 ( .A(n1071), .Y(n1063) );
  CLKBUFX2TS U150 ( .A(n1071), .Y(n1062) );
  CLKBUFX2TS U151 ( .A(n1075), .Y(n1046) );
  CLKBUFX2TS U152 ( .A(n1072), .Y(n1059) );
  CLKBUFX2TS U153 ( .A(n1072), .Y(n1058) );
  CLKBUFX2TS U154 ( .A(n1074), .Y(n1049) );
  CLKBUFX2TS U155 ( .A(n1074), .Y(n1050) );
  CLKBUFX2TS U156 ( .A(n1079), .Y(n1055) );
  CLKBUFX2TS U157 ( .A(n1073), .Y(n1053) );
  CLKBUFX2TS U158 ( .A(n1073), .Y(n1054) );
  CLKBUFX2TS U159 ( .A(n1080), .Y(n1069) );
  CLKBUFX2TS U160 ( .A(n1076), .Y(n1080) );
  CLKBUFX2TS U161 ( .A(n1078), .Y(n1075) );
  CLKBUFX2TS U162 ( .A(n1080), .Y(n1070) );
  INVX1TS U163 ( .A(n889), .Y(n890) );
  INVX1TS U164 ( .A(n691), .Y(n692) );
  INVX1TS U165 ( .A(n641), .Y(n642) );
  INVX1TS U166 ( .A(n951), .Y(n952) );
  INVX1TS U167 ( .A(n959), .Y(n960) );
  INVX1TS U168 ( .A(n703), .Y(n704) );
  INVX1TS U169 ( .A(n695), .Y(n696) );
  INVX1TS U170 ( .A(n949), .Y(n950) );
  INVX1TS U171 ( .A(n897), .Y(n898) );
  INVX1TS U172 ( .A(n737), .Y(n738) );
  INVX1TS U173 ( .A(n893), .Y(n894) );
  INVX1TS U174 ( .A(n699), .Y(n700) );
  INVX1TS U175 ( .A(n947), .Y(n948) );
  INVX1TS U176 ( .A(n1037), .Y(n1038) );
  INVX1TS U177 ( .A(n645), .Y(n646) );
  INVX1TS U178 ( .A(n967), .Y(n968) );
  INVX1TS U179 ( .A(n637), .Y(n638) );
  INVX1TS U180 ( .A(n971), .Y(n972) );
  INVX1TS U181 ( .A(n649), .Y(n650) );
  INVX1TS U182 ( .A(n711), .Y(n712) );
  INVX1TS U183 ( .A(n905), .Y(n906) );
  INVX1TS U184 ( .A(n911), .Y(n912) );
  INVX1TS U185 ( .A(n655), .Y(n656) );
  INVX1TS U186 ( .A(n715), .Y(n716) );
  INVX1TS U187 ( .A(n955), .Y(n956) );
  INVX1TS U188 ( .A(n653), .Y(n654) );
  INVX1TS U189 ( .A(n989), .Y(n990) );
  INVX1TS U190 ( .A(n915), .Y(n916) );
  INVX1TS U191 ( .A(n659), .Y(n660) );
  INVX1TS U192 ( .A(n697), .Y(n698) );
  INVX1TS U193 ( .A(n909), .Y(n910) );
  INVX1TS U194 ( .A(n919), .Y(n920) );
  INVX1TS U195 ( .A(n663), .Y(n664) );
  INVX1TS U196 ( .A(n593), .Y(n594) );
  INVX1TS U197 ( .A(n963), .Y(n964) );
  INVX1TS U198 ( .A(n707), .Y(n708) );
  INVX1TS U199 ( .A(n923), .Y(n924) );
  INVX1TS U200 ( .A(n901), .Y(n902) );
  INVX1TS U201 ( .A(n667), .Y(n668) );
  INVX1TS U202 ( .A(n849), .Y(n850) );
  INVX1TS U203 ( .A(n927), .Y(n928) );
  INVX1TS U204 ( .A(n671), .Y(n672) );
  INVX1TS U205 ( .A(n597), .Y(n598) );
  INVX1TS U206 ( .A(n853), .Y(n854) );
  INVX1TS U207 ( .A(n931), .Y(n932) );
  INVX1TS U208 ( .A(n675), .Y(n676) );
  INVX1TS U209 ( .A(n601), .Y(n602) );
  INVX1TS U210 ( .A(n935), .Y(n936) );
  INVX1TS U211 ( .A(n733), .Y(n734) );
  INVX1TS U212 ( .A(n679), .Y(n680) );
  INVX1TS U213 ( .A(n953), .Y(n954) );
  INVX1TS U214 ( .A(n857), .Y(n858) );
  INVX1TS U215 ( .A(n939), .Y(n940) );
  INVX1TS U216 ( .A(n683), .Y(n684) );
  INVX1TS U217 ( .A(n879), .Y(n880) );
  INVX1TS U218 ( .A(n605), .Y(n606) );
  INVX1TS U219 ( .A(n623), .Y(n624) );
  INVX1TS U220 ( .A(n883), .Y(n884) );
  INVX1TS U221 ( .A(n861), .Y(n862) );
  INVX1TS U222 ( .A(n627), .Y(n628) );
  INVX1TS U223 ( .A(n609), .Y(n610) );
  INVX1TS U224 ( .A(n887), .Y(n888) );
  INVX1TS U225 ( .A(n631), .Y(n632) );
  INVX1TS U226 ( .A(n701), .Y(n702) );
  INVX1TS U227 ( .A(n865), .Y(n866) );
  INVX1TS U228 ( .A(n891), .Y(n892) );
  INVX1TS U229 ( .A(n635), .Y(n636) );
  INVX1TS U230 ( .A(n895), .Y(n896) );
  INVX1TS U231 ( .A(n613), .Y(n614) );
  INVX1TS U232 ( .A(n639), .Y(n640) );
  INVX1TS U233 ( .A(n985), .Y(n986) );
  INVX1TS U234 ( .A(n899), .Y(n900) );
  INVX1TS U235 ( .A(n869), .Y(n870) );
  INVX1TS U236 ( .A(n643), .Y(n644) );
  INVX1TS U237 ( .A(n903), .Y(n904) );
  INVX1TS U238 ( .A(n957), .Y(n958) );
  INVX1TS U239 ( .A(n647), .Y(n648) );
  INVX1TS U240 ( .A(n617), .Y(n618) );
  INVX1TS U241 ( .A(n907), .Y(n908) );
  INVX1TS U242 ( .A(n651), .Y(n652) );
  INVX1TS U243 ( .A(n873), .Y(n874) );
  INVX1TS U244 ( .A(n721), .Y(n722) );
  INVX1TS U245 ( .A(n847), .Y(n848) );
  INVX1TS U246 ( .A(n621), .Y(n622) );
  INVX1TS U247 ( .A(n591), .Y(n592) );
  INVX1TS U248 ( .A(n781), .Y(n782) );
  INVX1TS U249 ( .A(n705), .Y(n706) );
  INVX1TS U250 ( .A(n1001), .Y(n1002) );
  INVX1TS U251 ( .A(n961), .Y(n962) );
  INVX1TS U252 ( .A(n1033), .Y(n1034) );
  INVX1TS U253 ( .A(n777), .Y(n778) );
  INVX1TS U254 ( .A(n709), .Y(n710) );
  INVX1TS U255 ( .A(n965), .Y(n966) );
  INVX1TS U256 ( .A(n1029), .Y(n1030) );
  INVX1TS U257 ( .A(n773), .Y(n774) );
  INVX1TS U258 ( .A(n1025), .Y(n1026) );
  INVX1TS U259 ( .A(n713), .Y(n714) );
  INVX1TS U260 ( .A(n769), .Y(n770) );
  INVX1TS U261 ( .A(n745), .Y(n746) );
  INVX1TS U262 ( .A(n1021), .Y(n1022) );
  INVX1TS U263 ( .A(n969), .Y(n970) );
  INVX1TS U264 ( .A(n765), .Y(n766) );
  INVX1TS U265 ( .A(n717), .Y(n718) );
  INVX1TS U266 ( .A(n1017), .Y(n1018) );
  INVX1TS U267 ( .A(n761), .Y(n762) );
  INVX1TS U268 ( .A(n749), .Y(n750) );
  INVX1TS U269 ( .A(n973), .Y(n974) );
  INVX1TS U270 ( .A(n1013), .Y(n1014) );
  INVX1TS U271 ( .A(n757), .Y(n758) );
  INVX1TS U272 ( .A(n657), .Y(n658) );
  INVX1TS U273 ( .A(n1009), .Y(n1010) );
  INVX1TS U274 ( .A(n753), .Y(n754) );
  INVX1TS U275 ( .A(n913), .Y(n914) );
  INVX1TS U276 ( .A(n1007), .Y(n1008) );
  INVX1TS U277 ( .A(n751), .Y(n752) );
  INVX1TS U278 ( .A(n661), .Y(n662) );
  INVX1TS U279 ( .A(n917), .Y(n918) );
  INVX1TS U280 ( .A(n1011), .Y(n1012) );
  INVX1TS U281 ( .A(n755), .Y(n756) );
  INVX1TS U282 ( .A(n665), .Y(n666) );
  INVX1TS U283 ( .A(n997), .Y(n998) );
  INVX1TS U284 ( .A(n1005), .Y(n1006) );
  INVX1TS U285 ( .A(n1015), .Y(n1016) );
  INVX1TS U286 ( .A(n759), .Y(n760) );
  INVX1TS U287 ( .A(n921), .Y(n922) );
  INVX1TS U288 ( .A(n1019), .Y(n1020) );
  INVX1TS U289 ( .A(n763), .Y(n764) );
  INVX1TS U290 ( .A(n669), .Y(n670) );
  INVX1TS U291 ( .A(n1023), .Y(n1024) );
  INVX1TS U292 ( .A(n767), .Y(n768) );
  INVX1TS U293 ( .A(n925), .Y(n926) );
  INVX1TS U294 ( .A(n1027), .Y(n1028) );
  INVX1TS U295 ( .A(n771), .Y(n772) );
  INVX1TS U296 ( .A(n673), .Y(n674) );
  INVX1TS U297 ( .A(n1031), .Y(n1032) );
  INVX1TS U298 ( .A(n775), .Y(n776) );
  INVX1TS U299 ( .A(n929), .Y(n930) );
  INVX1TS U300 ( .A(n1035), .Y(n1036) );
  INVX1TS U301 ( .A(n779), .Y(n780) );
  INVX1TS U302 ( .A(n741), .Y(n742) );
  INVX1TS U303 ( .A(n689), .Y(n690) );
  INVX1TS U304 ( .A(n677), .Y(n678) );
  INVX1TS U305 ( .A(n975), .Y(n976) );
  INVX1TS U306 ( .A(n719), .Y(n720) );
  INVX1TS U307 ( .A(n933), .Y(n934) );
  INVX1TS U308 ( .A(n681), .Y(n682) );
  INVX1TS U309 ( .A(n979), .Y(n980) );
  INVX1TS U310 ( .A(n723), .Y(n724) );
  INVX1TS U311 ( .A(n937), .Y(n938) );
  INVX1TS U312 ( .A(n983), .Y(n984) );
  INVX1TS U313 ( .A(n727), .Y(n728) );
  INVX1TS U314 ( .A(n685), .Y(n686) );
  INVX1TS U315 ( .A(n987), .Y(n988) );
  INVX1TS U316 ( .A(n731), .Y(n732) );
  INVX1TS U317 ( .A(n945), .Y(n946) );
  INVX1TS U318 ( .A(n941), .Y(n942) );
  INVX1TS U319 ( .A(n991), .Y(n992) );
  INVX1TS U320 ( .A(n735), .Y(n736) );
  INVX1TS U321 ( .A(n625), .Y(n626) );
  INVX1TS U322 ( .A(n881), .Y(n882) );
  INVX1TS U323 ( .A(n995), .Y(n996) );
  INVX1TS U324 ( .A(n739), .Y(n740) );
  INVX1TS U325 ( .A(n993), .Y(n994) );
  INVX1TS U326 ( .A(n999), .Y(n1000) );
  INVX1TS U327 ( .A(n629), .Y(n630) );
  INVX1TS U328 ( .A(n743), .Y(n744) );
  INVX1TS U329 ( .A(n1003), .Y(n1004) );
  INVX1TS U330 ( .A(n885), .Y(n886) );
  INVX1TS U331 ( .A(n747), .Y(n748) );
  INVX1TS U332 ( .A(n633), .Y(n634) );
  INVX1TS U333 ( .A(n943), .Y(n944) );
  INVX1TS U334 ( .A(n693), .Y(n694) );
  INVX1TS U335 ( .A(n687), .Y(n688) );
  INVX1TS U336 ( .A(n789), .Y(n790) );
  INVX1TS U337 ( .A(n607), .Y(n608) );
  INVX1TS U338 ( .A(n803), .Y(n804) );
  INVX1TS U339 ( .A(n725), .Y(n726) );
  INVX1TS U340 ( .A(n543), .Y(n544) );
  INVX1TS U341 ( .A(n587), .Y(n588) );
  INVX1TS U342 ( .A(n565), .Y(n566) );
  INVX1TS U343 ( .A(n863), .Y(n864) );
  INVX1TS U344 ( .A(n547), .Y(n548) );
  INVX1TS U345 ( .A(n585), .Y(n586) );
  INVX1TS U346 ( .A(n977), .Y(n978) );
  INVX1TS U347 ( .A(n583), .Y(n584) );
  INVX1TS U348 ( .A(n537), .Y(n538) );
  INVX1TS U349 ( .A(n815), .Y(n816) );
  INVX1TS U350 ( .A(n841), .Y(n842) );
  INVX1TS U351 ( .A(n533), .Y(n534) );
  INVX1TS U352 ( .A(n573), .Y(n574) );
  INVX1TS U353 ( .A(n839), .Y(n840) );
  INVX1TS U354 ( .A(n807), .Y(n808) );
  INVX1TS U355 ( .A(n799), .Y(n800) );
  INVX1TS U356 ( .A(n825), .Y(n826) );
  INVX1TS U357 ( .A(n603), .Y(n604) );
  INVX1TS U358 ( .A(n551), .Y(n552) );
  INVX1TS U359 ( .A(n559), .Y(n560) );
  INVX1TS U360 ( .A(n793), .Y(n794) );
  INVX1TS U361 ( .A(n867), .Y(n868) );
  INVX1TS U362 ( .A(n821), .Y(n822) );
  INVX1TS U363 ( .A(n619), .Y(n620) );
  INVX1TS U364 ( .A(n811), .Y(n812) );
  INVX1TS U365 ( .A(n579), .Y(n580) );
  INVX1TS U366 ( .A(n859), .Y(n860) );
  INVX1TS U367 ( .A(n837), .Y(n838) );
  INVX1TS U368 ( .A(n539), .Y(n540) );
  INVX1TS U369 ( .A(n555), .Y(n556) );
  INVX1TS U370 ( .A(n835), .Y(n836) );
  INVX1TS U371 ( .A(n783), .Y(n784) );
  INVX1TS U372 ( .A(n589), .Y(n590) );
  INVX1TS U373 ( .A(n817), .Y(n818) );
  INVX1TS U374 ( .A(n729), .Y(n730) );
  INVX1TS U375 ( .A(n611), .Y(n612) );
  INVX1TS U376 ( .A(n599), .Y(n600) );
  INVX1TS U377 ( .A(n813), .Y(n814) );
  INVX1TS U378 ( .A(n541), .Y(n542) );
  INVX1TS U379 ( .A(n795), .Y(n796) );
  INVX1TS U380 ( .A(n819), .Y(n820) );
  INVX1TS U381 ( .A(n875), .Y(n876) );
  INVX1TS U382 ( .A(n843), .Y(n844) );
  INVX1TS U383 ( .A(n829), .Y(n830) );
  INVX1TS U384 ( .A(n575), .Y(n576) );
  INVX1TS U385 ( .A(n557), .Y(n558) );
  INVX1TS U386 ( .A(n527), .Y(n528) );
  INVX1TS U387 ( .A(n615), .Y(n616) );
  INVX1TS U388 ( .A(n785), .Y(n786) );
  INVX1TS U389 ( .A(n981), .Y(n982) );
  INVX1TS U390 ( .A(n577), .Y(n578) );
  INVX1TS U391 ( .A(n833), .Y(n834) );
  INVX1TS U392 ( .A(n855), .Y(n856) );
  INVX1TS U393 ( .A(n595), .Y(n596) );
  INVX1TS U394 ( .A(n561), .Y(n562) );
  INVX1TS U395 ( .A(n581), .Y(n582) );
  INVX1TS U396 ( .A(n831), .Y(n832) );
  INVX1TS U397 ( .A(n827), .Y(n828) );
  INVX1TS U398 ( .A(n553), .Y(n554) );
  INVX1TS U399 ( .A(n809), .Y(n810) );
  INVX1TS U400 ( .A(n797), .Y(n798) );
  INVX1TS U401 ( .A(n563), .Y(n564) );
  INVX1TS U402 ( .A(n569), .Y(n570) );
  INVX1TS U403 ( .A(n877), .Y(n878) );
  INVX1TS U404 ( .A(n845), .Y(n846) );
  INVX1TS U405 ( .A(n535), .Y(n536) );
  INVX1TS U406 ( .A(n529), .Y(n530) );
  INVX1TS U407 ( .A(n567), .Y(n568) );
  INVX1TS U408 ( .A(n823), .Y(n824) );
  INVX1TS U409 ( .A(n791), .Y(n792) );
  INVX1TS U410 ( .A(n805), .Y(n806) );
  INVX1TS U411 ( .A(n787), .Y(n788) );
  INVX1TS U412 ( .A(n571), .Y(n572) );
  INVX1TS U413 ( .A(n545), .Y(n546) );
  INVX1TS U414 ( .A(n871), .Y(n872) );
  INVX1TS U415 ( .A(n549), .Y(n550) );
  INVX1TS U416 ( .A(n851), .Y(n852) );
  INVX1TS U417 ( .A(n531), .Y(n532) );
  INVX1TS U418 ( .A(n801), .Y(n802) );
  INVXLTS U419 ( .A(\ux33/n10 ), .Y(n525) );
  INVXLTS U420 ( .A(n525), .Y(n526) );
  INVXLTS U421 ( .A(text_in_r[64]), .Y(n527) );
  INVXLTS U422 ( .A(text_in_r[63]), .Y(n529) );
  INVXLTS U423 ( .A(text_in_r[65]), .Y(n531) );
  INVXLTS U424 ( .A(text_in_r[62]), .Y(n533) );
  INVXLTS U425 ( .A(text_in_r[66]), .Y(n535) );
  INVXLTS U426 ( .A(text_in_r[61]), .Y(n537) );
  INVXLTS U427 ( .A(text_in_r[67]), .Y(n539) );
  INVXLTS U428 ( .A(text_in_r[60]), .Y(n541) );
  INVXLTS U429 ( .A(text_in_r[68]), .Y(n543) );
  INVXLTS U430 ( .A(text_in_r[59]), .Y(n545) );
  INVXLTS U431 ( .A(text_in_r[69]), .Y(n547) );
  INVXLTS U432 ( .A(text_in_r[58]), .Y(n549) );
  INVXLTS U433 ( .A(text_in_r[70]), .Y(n551) );
  INVXLTS U434 ( .A(text_in_r[57]), .Y(n553) );
  INVXLTS U435 ( .A(text_in_r[71]), .Y(n555) );
  INVXLTS U436 ( .A(text_in_r[56]), .Y(n557) );
  INVXLTS U437 ( .A(text_in_r[72]), .Y(n559) );
  INVXLTS U438 ( .A(text_in_r[55]), .Y(n561) );
  INVXLTS U439 ( .A(text_in_r[73]), .Y(n563) );
  INVXLTS U440 ( .A(text_in_r[54]), .Y(n565) );
  INVXLTS U441 ( .A(text_in_r[74]), .Y(n567) );
  INVXLTS U442 ( .A(text_in_r[53]), .Y(n569) );
  INVXLTS U443 ( .A(text_in_r[75]), .Y(n571) );
  INVXLTS U444 ( .A(text_in_r[52]), .Y(n573) );
  INVXLTS U445 ( .A(text_in_r[76]), .Y(n575) );
  INVXLTS U446 ( .A(text_in_r[51]), .Y(n577) );
  INVXLTS U447 ( .A(text_in_r[77]), .Y(n579) );
  INVXLTS U448 ( .A(text_in_r[50]), .Y(n581) );
  INVXLTS U449 ( .A(text_in_r[78]), .Y(n583) );
  INVXLTS U450 ( .A(text_in_r[49]), .Y(n585) );
  INVXLTS U451 ( .A(text_in_r[79]), .Y(n587) );
  INVXLTS U452 ( .A(text_in_r[48]), .Y(n589) );
  INVXLTS U453 ( .A(text_in_r[80]), .Y(n591) );
  INVXLTS U454 ( .A(text_in_r[47]), .Y(n593) );
  INVXLTS U455 ( .A(text_in_r[81]), .Y(n595) );
  INVXLTS U456 ( .A(text_in_r[46]), .Y(n597) );
  INVXLTS U457 ( .A(text_in_r[82]), .Y(n599) );
  INVXLTS U458 ( .A(text_in_r[45]), .Y(n601) );
  INVXLTS U459 ( .A(text_in_r[83]), .Y(n603) );
  INVXLTS U460 ( .A(text_in_r[44]), .Y(n605) );
  INVXLTS U461 ( .A(text_in_r[84]), .Y(n607) );
  INVXLTS U462 ( .A(text_in_r[43]), .Y(n609) );
  INVXLTS U463 ( .A(text_in_r[85]), .Y(n611) );
  INVXLTS U464 ( .A(text_in_r[42]), .Y(n613) );
  INVXLTS U465 ( .A(text_in_r[86]), .Y(n615) );
  INVXLTS U466 ( .A(text_in_r[41]), .Y(n617) );
  INVXLTS U467 ( .A(text_in_r[87]), .Y(n619) );
  INVXLTS U468 ( .A(text_in_r[40]), .Y(n621) );
  INVXLTS U469 ( .A(text_in_r[88]), .Y(n623) );
  INVXLTS U470 ( .A(text_in_r[39]), .Y(n625) );
  INVXLTS U471 ( .A(text_in_r[89]), .Y(n627) );
  INVXLTS U472 ( .A(text_in_r[38]), .Y(n629) );
  INVXLTS U473 ( .A(text_in_r[90]), .Y(n631) );
  INVXLTS U474 ( .A(text_in_r[37]), .Y(n633) );
  INVXLTS U475 ( .A(text_in_r[91]), .Y(n635) );
  INVXLTS U476 ( .A(text_in_r[36]), .Y(n637) );
  INVXLTS U477 ( .A(text_in_r[92]), .Y(n639) );
  INVXLTS U478 ( .A(text_in_r[35]), .Y(n641) );
  INVXLTS U479 ( .A(text_in_r[93]), .Y(n643) );
  INVXLTS U480 ( .A(text_in_r[34]), .Y(n645) );
  INVXLTS U481 ( .A(text_in_r[94]), .Y(n647) );
  INVXLTS U482 ( .A(text_in_r[33]), .Y(n649) );
  INVXLTS U483 ( .A(text_in_r[95]), .Y(n651) );
  INVXLTS U484 ( .A(text_in_r[32]), .Y(n653) );
  INVXLTS U485 ( .A(text_in_r[96]), .Y(n655) );
  INVXLTS U486 ( .A(text_in_r[31]), .Y(n657) );
  INVXLTS U487 ( .A(text_in_r[97]), .Y(n659) );
  INVXLTS U488 ( .A(text_in_r[30]), .Y(n661) );
  INVXLTS U489 ( .A(text_in_r[98]), .Y(n663) );
  INVXLTS U490 ( .A(text_in_r[29]), .Y(n665) );
  INVXLTS U491 ( .A(text_in_r[99]), .Y(n667) );
  INVXLTS U492 ( .A(text_in_r[28]), .Y(n669) );
  INVXLTS U493 ( .A(text_in_r[100]), .Y(n671) );
  INVXLTS U494 ( .A(text_in_r[27]), .Y(n673) );
  INVXLTS U495 ( .A(text_in_r[101]), .Y(n675) );
  INVXLTS U496 ( .A(text_in_r[26]), .Y(n677) );
  INVXLTS U497 ( .A(text_in_r[102]), .Y(n679) );
  INVXLTS U498 ( .A(text_in_r[25]), .Y(n681) );
  INVXLTS U499 ( .A(text_in_r[103]), .Y(n683) );
  INVXLTS U500 ( .A(text_in_r[24]), .Y(n685) );
  INVXLTS U501 ( .A(text_in_r[104]), .Y(n687) );
  INVXLTS U502 ( .A(text_in_r[23]), .Y(n689) );
  INVXLTS U503 ( .A(text_in_r[105]), .Y(n691) );
  INVXLTS U504 ( .A(text_in_r[22]), .Y(n693) );
  INVXLTS U505 ( .A(text_in_r[106]), .Y(n695) );
  INVXLTS U506 ( .A(text_in_r[21]), .Y(n697) );
  INVXLTS U507 ( .A(text_in_r[107]), .Y(n699) );
  INVXLTS U508 ( .A(text_in_r[20]), .Y(n701) );
  INVXLTS U509 ( .A(text_in_r[108]), .Y(n703) );
  INVXLTS U510 ( .A(text_in_r[19]), .Y(n705) );
  INVXLTS U511 ( .A(text_in_r[109]), .Y(n707) );
  INVXLTS U512 ( .A(text_in_r[18]), .Y(n709) );
  INVXLTS U513 ( .A(text_in_r[110]), .Y(n711) );
  INVXLTS U514 ( .A(text_in_r[17]), .Y(n713) );
  INVXLTS U515 ( .A(text_in_r[111]), .Y(n715) );
  INVXLTS U516 ( .A(text_in_r[16]), .Y(n717) );
  INVXLTS U517 ( .A(text_in_r[112]), .Y(n719) );
  INVXLTS U518 ( .A(text_in_r[15]), .Y(n721) );
  INVXLTS U519 ( .A(text_in_r[113]), .Y(n723) );
  INVXLTS U520 ( .A(text_in_r[14]), .Y(n725) );
  INVXLTS U521 ( .A(text_in_r[114]), .Y(n727) );
  INVXLTS U522 ( .A(text_in_r[13]), .Y(n729) );
  INVXLTS U523 ( .A(text_in_r[115]), .Y(n731) );
  INVXLTS U524 ( .A(text_in_r[12]), .Y(n733) );
  INVXLTS U525 ( .A(text_in_r[116]), .Y(n735) );
  INVXLTS U526 ( .A(text_in_r[11]), .Y(n737) );
  INVXLTS U527 ( .A(text_in_r[117]), .Y(n739) );
  INVXLTS U528 ( .A(text_in_r[10]), .Y(n741) );
  INVXLTS U529 ( .A(text_in_r[118]), .Y(n743) );
  INVXLTS U530 ( .A(text_in_r[9]), .Y(n745) );
  INVXLTS U531 ( .A(text_in_r[119]), .Y(n747) );
  INVXLTS U532 ( .A(text_in_r[8]), .Y(n749) );
  INVXLTS U533 ( .A(text_in_r[120]), .Y(n751) );
  INVXLTS U534 ( .A(text_in_r[7]), .Y(n753) );
  INVXLTS U535 ( .A(text_in_r[121]), .Y(n755) );
  INVXLTS U536 ( .A(text_in_r[6]), .Y(n757) );
  INVXLTS U537 ( .A(text_in_r[122]), .Y(n759) );
  INVXLTS U538 ( .A(text_in_r[5]), .Y(n761) );
  INVXLTS U539 ( .A(text_in_r[123]), .Y(n763) );
  INVXLTS U540 ( .A(text_in_r[4]), .Y(n765) );
  INVXLTS U541 ( .A(text_in_r[124]), .Y(n767) );
  INVXLTS U542 ( .A(text_in_r[3]), .Y(n769) );
  INVXLTS U543 ( .A(text_in_r[125]), .Y(n771) );
  INVXLTS U544 ( .A(text_in_r[2]), .Y(n773) );
  INVXLTS U545 ( .A(text_in_r[126]), .Y(n775) );
  INVXLTS U546 ( .A(text_in_r[1]), .Y(n777) );
  INVXLTS U547 ( .A(text_in_r[127]), .Y(n779) );
  INVXLTS U548 ( .A(text_in_r[0]), .Y(n781) );
  INVXLTS U549 ( .A(w1[0]), .Y(n783) );
  INVXLTS U550 ( .A(w2[31]), .Y(n785) );
  INVXLTS U551 ( .A(w1[1]), .Y(n787) );
  INVXLTS U552 ( .A(w2[30]), .Y(n789) );
  INVXLTS U553 ( .A(w1[2]), .Y(n791) );
  INVXLTS U554 ( .A(w2[29]), .Y(n793) );
  INVXLTS U555 ( .A(w1[3]), .Y(n795) );
  INVXLTS U556 ( .A(w2[28]), .Y(n797) );
  INVXLTS U557 ( .A(w1[4]), .Y(n799) );
  INVXLTS U558 ( .A(w2[27]), .Y(n801) );
  INVXLTS U559 ( .A(w1[5]), .Y(n803) );
  INVXLTS U560 ( .A(w2[26]), .Y(n805) );
  INVXLTS U561 ( .A(w1[6]), .Y(n807) );
  INVXLTS U562 ( .A(w2[25]), .Y(n809) );
  INVXLTS U563 ( .A(w1[7]), .Y(n811) );
  INVXLTS U564 ( .A(w2[24]), .Y(n813) );
  INVXLTS U565 ( .A(w1[8]), .Y(n815) );
  INVXLTS U566 ( .A(w2[23]), .Y(n817) );
  INVXLTS U567 ( .A(w1[9]), .Y(n819) );
  INVXLTS U568 ( .A(w2[22]), .Y(n821) );
  INVXLTS U569 ( .A(w1[10]), .Y(n823) );
  INVXLTS U570 ( .A(w2[21]), .Y(n825) );
  INVXLTS U571 ( .A(w1[11]), .Y(n827) );
  INVXLTS U572 ( .A(w2[20]), .Y(n829) );
  INVXLTS U573 ( .A(w1[12]), .Y(n831) );
  INVXLTS U574 ( .A(w2[19]), .Y(n833) );
  INVXLTS U575 ( .A(w1[13]), .Y(n835) );
  INVXLTS U576 ( .A(w2[18]), .Y(n837) );
  INVXLTS U577 ( .A(w1[14]), .Y(n839) );
  INVXLTS U578 ( .A(w2[17]), .Y(n841) );
  INVXLTS U579 ( .A(w1[15]), .Y(n843) );
  INVXLTS U580 ( .A(w2[16]), .Y(n845) );
  INVXLTS U581 ( .A(w1[16]), .Y(n847) );
  INVXLTS U582 ( .A(w2[15]), .Y(n849) );
  INVXLTS U583 ( .A(w1[17]), .Y(n851) );
  INVXLTS U584 ( .A(w2[14]), .Y(n853) );
  INVXLTS U585 ( .A(w1[18]), .Y(n855) );
  INVXLTS U586 ( .A(w2[13]), .Y(n857) );
  INVXLTS U587 ( .A(w1[19]), .Y(n859) );
  INVXLTS U588 ( .A(w2[12]), .Y(n861) );
  INVXLTS U589 ( .A(w1[20]), .Y(n863) );
  INVXLTS U590 ( .A(w2[11]), .Y(n865) );
  INVXLTS U591 ( .A(w1[21]), .Y(n867) );
  INVXLTS U592 ( .A(w2[10]), .Y(n869) );
  INVXLTS U593 ( .A(w1[22]), .Y(n871) );
  INVXLTS U594 ( .A(w2[9]), .Y(n873) );
  INVXLTS U595 ( .A(w1[23]), .Y(n875) );
  INVXLTS U596 ( .A(w2[8]), .Y(n877) );
  INVXLTS U597 ( .A(w1[24]), .Y(n879) );
  INVXLTS U598 ( .A(w2[7]), .Y(n881) );
  INVXLTS U599 ( .A(w1[25]), .Y(n883) );
  INVXLTS U600 ( .A(w2[6]), .Y(n885) );
  INVXLTS U601 ( .A(w1[26]), .Y(n887) );
  INVXLTS U602 ( .A(w2[5]), .Y(n889) );
  INVXLTS U603 ( .A(w1[27]), .Y(n891) );
  INVXLTS U604 ( .A(w2[4]), .Y(n893) );
  INVXLTS U605 ( .A(w1[28]), .Y(n895) );
  INVXLTS U606 ( .A(w2[3]), .Y(n897) );
  INVXLTS U607 ( .A(w1[29]), .Y(n899) );
  INVXLTS U608 ( .A(w2[2]), .Y(n901) );
  INVXLTS U609 ( .A(w1[30]), .Y(n903) );
  INVXLTS U610 ( .A(w2[1]), .Y(n905) );
  INVXLTS U611 ( .A(w1[31]), .Y(n907) );
  INVXLTS U612 ( .A(w2[0]), .Y(n909) );
  INVXLTS U613 ( .A(w0[0]), .Y(n911) );
  INVXLTS U614 ( .A(w3[31]), .Y(n913) );
  INVXLTS U615 ( .A(w0[1]), .Y(n915) );
  INVXLTS U616 ( .A(w3[30]), .Y(n917) );
  INVXLTS U617 ( .A(w0[2]), .Y(n919) );
  INVXLTS U618 ( .A(w3[29]), .Y(n921) );
  INVXLTS U619 ( .A(w0[3]), .Y(n923) );
  INVXLTS U620 ( .A(w3[28]), .Y(n925) );
  INVXLTS U621 ( .A(w0[4]), .Y(n927) );
  INVXLTS U622 ( .A(w3[27]), .Y(n929) );
  INVXLTS U623 ( .A(w0[5]), .Y(n931) );
  INVXLTS U624 ( .A(w3[26]), .Y(n933) );
  INVXLTS U625 ( .A(w0[6]), .Y(n935) );
  INVXLTS U626 ( .A(w3[25]), .Y(n937) );
  INVXLTS U627 ( .A(w0[7]), .Y(n939) );
  INVXLTS U628 ( .A(w3[24]), .Y(n941) );
  INVXLTS U629 ( .A(w0[8]), .Y(n943) );
  INVXLTS U630 ( .A(w3[23]), .Y(n945) );
  INVXLTS U631 ( .A(w0[9]), .Y(n947) );
  INVXLTS U632 ( .A(w3[22]), .Y(n949) );
  INVXLTS U633 ( .A(w0[10]), .Y(n951) );
  INVXLTS U634 ( .A(w3[21]), .Y(n953) );
  INVXLTS U635 ( .A(w0[11]), .Y(n955) );
  INVXLTS U636 ( .A(w3[20]), .Y(n957) );
  INVXLTS U637 ( .A(w0[12]), .Y(n959) );
  INVXLTS U638 ( .A(w3[19]), .Y(n961) );
  INVXLTS U639 ( .A(w0[13]), .Y(n963) );
  INVXLTS U640 ( .A(w3[18]), .Y(n965) );
  INVXLTS U641 ( .A(w0[14]), .Y(n967) );
  INVXLTS U642 ( .A(w3[17]), .Y(n969) );
  INVXLTS U643 ( .A(w0[15]), .Y(n971) );
  INVXLTS U644 ( .A(w3[16]), .Y(n973) );
  INVXLTS U645 ( .A(w0[16]), .Y(n975) );
  INVXLTS U646 ( .A(w3[15]), .Y(n977) );
  INVXLTS U647 ( .A(w0[17]), .Y(n979) );
  INVXLTS U648 ( .A(w3[14]), .Y(n981) );
  INVXLTS U649 ( .A(w0[18]), .Y(n983) );
  INVXLTS U650 ( .A(w3[13]), .Y(n985) );
  INVXLTS U651 ( .A(w0[19]), .Y(n987) );
  INVXLTS U652 ( .A(w3[12]), .Y(n989) );
  INVXLTS U653 ( .A(w0[20]), .Y(n991) );
  INVXLTS U654 ( .A(w3[11]), .Y(n993) );
  INVXLTS U655 ( .A(w0[21]), .Y(n995) );
  INVXLTS U656 ( .A(w3[10]), .Y(n997) );
  INVXLTS U657 ( .A(w0[22]), .Y(n999) );
  INVXLTS U658 ( .A(w3[9]), .Y(n1001) );
  INVXLTS U659 ( .A(w0[23]), .Y(n1003) );
  INVXLTS U660 ( .A(w3[8]), .Y(n1005) );
  INVXLTS U661 ( .A(w0[24]), .Y(n1007) );
  INVXLTS U662 ( .A(w3[7]), .Y(n1009) );
  INVXLTS U663 ( .A(w0[25]), .Y(n1011) );
  INVXLTS U664 ( .A(w3[6]), .Y(n1013) );
  INVXLTS U665 ( .A(w0[26]), .Y(n1015) );
  INVXLTS U666 ( .A(w3[5]), .Y(n1017) );
  INVXLTS U667 ( .A(w0[27]), .Y(n1019) );
  INVXLTS U668 ( .A(w3[4]), .Y(n1021) );
  INVXLTS U669 ( .A(w0[28]), .Y(n1023) );
  INVXLTS U670 ( .A(w3[3]), .Y(n1025) );
  INVXLTS U671 ( .A(w0[29]), .Y(n1027) );
  INVXLTS U672 ( .A(w3[2]), .Y(n1029) );
  INVXLTS U673 ( .A(w0[30]), .Y(n1031) );
  INVXLTS U674 ( .A(w3[1]), .Y(n1033) );
  INVXLTS U675 ( .A(w0[31]), .Y(n1035) );
  INVXLTS U676 ( .A(w3[0]), .Y(n1037) );
  CLKBUFX2TS U677 ( .A(n526), .Y(n1079) );
  CLKBUFX2TS U678 ( .A(n526), .Y(n1077) );
  CLKBUFX2TS U679 ( .A(n526), .Y(n1076) );
  CLKBUFX2TS U680 ( .A(n1077), .Y(n1045) );
  CLKBUFX2TS U681 ( .A(n1077), .Y(n1039) );
  CLKBUFX2TS U682 ( .A(n1076), .Y(n1042) );
  CLKBUFX2TS U683 ( .A(n1076), .Y(n1040) );
  CLKBUFX2TS U684 ( .A(n1076), .Y(n1041) );
endmodule

