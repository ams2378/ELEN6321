.TEMP 25
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2

xu8 clk d_bar_o qbar_o DFFQX1TS
.END
