library verilog;
use verilog.vl_types.all;
entity wddl_dflipflop_tb is
end wddl_dflipflop_tb;
