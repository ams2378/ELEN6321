.subckt aes_xor sa_i7 sa_i6 sa_i5 sa_i4 sa_i3 sa_i2 sa_i1 sa_i0 
+ sa_o7 sa_o6 sa_o5 sa_o4 sa_o3 sa_o2 sa_o1 sa_o0 
+ text_in7 text_in6 text_in5 text_in4 text_in3 text_in2 text_in1 text_in0 
+ w_i7 w_i6 w_i5 w_i4 w_i3 w_i2 w_i1 w_i0 clk ld_r gnd vdd
x1XOR2X1TS n8 n102 n86 gnd vdd XOR2X1TS
x2XOR2X1TS n7 n98 n82 gnd vdd XOR2X1TS
x3XOR2X1TS n6 n94 n78 gnd vdd XOR2X1TS
x4XOR2X1TS n2 n108 n92 gnd vdd XOR2X1TS
x5XOR2X1TS n5 n96 n80 gnd vdd XOR2X1TS
x6XOR2X1TS n4 n100 n84 gnd vdd XOR2X1TS
x7XOR2X1TS n3 n104 n88 gnd vdd XOR2X1TS
x8XOR2X1TS n9 n106 n90 gnd vdd XOR2X1TS
x9SDFFQXLTS sa_o7 clk sa_i7 n110 n2 gnd vdd SDFFQXLTS
x10SDFFQXLTS sa_o6 clk sa_i6 n111 n3 gnd vdd SDFFQXLTS
x11SDFFQXLTS sa_o5 clk sa_i5 n111 n4 gnd vdd SDFFQXLTS
x12SDFFQXLTS sa_o4 clk sa_i4 n110 n5 gnd vdd SDFFQXLTS
x13SDFFQXLTS sa_o3 clk sa_i3 n111 n6 gnd vdd SDFFQXLTS
x14SDFFQXLTS sa_o2 clk sa_i2 n110 n7 gnd vdd SDFFQXLTS
x15SDFFQXLTS sa_o1 clk sa_i1 n110 n8 gnd vdd SDFFQXLTS
x16SDFFQXLTS sa_o0 clk sa_i0 n111 n9 gnd vdd SDFFQXLTS
x17INVX1TS n92 n91 gnd vdd INVX1TS
x18INVX1TS n88 n87 gnd vdd INVX1TS
x19INVX1TS n100 n99 gnd vdd INVX1TS
x20INVX1TS n84 n83 gnd vdd INVX1TS
x21INVX1TS n96 n95 gnd vdd INVX1TS
x22INVX1TS n111 n109 gnd vdd INVX1TS
x23INVX1TS n108 n107 gnd vdd INVX1TS
x24INVX1TS n80 n79 gnd vdd INVX1TS
x25INVX1TS n104 n103 gnd vdd INVX1TS
x26INVX1TS n110 n109 gnd vdd INVX1TS
x27INVX1TS n102 n101 gnd vdd INVX1TS
x28INVX1TS n86 n85 gnd vdd INVX1TS
x29INVX1TS n90 n89 gnd vdd INVX1TS
x30INVX1TS n98 n97 gnd vdd INVX1TS
x31INVX1TS n106 n105 gnd vdd INVX1TS
x32INVX1TS n82 n81 gnd vdd INVX1TS
x33INVX1TS n94 n93 gnd vdd INVX1TS
x34INVX1TS n78 n77 gnd vdd INVX1TS
x35INVXLTS n77 text_in3 gnd vdd INVXLTS
x36INVXLTS n79 text_in4 gnd vdd INVXLTS
x37INVXLTS n81 text_in2 gnd vdd INVXLTS
x38INVXLTS n83 text_in5 gnd vdd INVXLTS
x39INVXLTS n85 text_in1 gnd vdd INVXLTS
x40INVXLTS n87 text_in6 gnd vdd INVXLTS
x41INVXLTS n89 text_in0 gnd vdd INVXLTS
x42INVXLTS n91 text_in7 gnd vdd INVXLTS
x43INVXLTS n93 w_i3 gnd vdd INVXLTS
x44INVXLTS n95 w_i4 gnd vdd INVXLTS
x45INVXLTS n97 w_i2 gnd vdd INVXLTS
x46INVXLTS n99 w_i5 gnd vdd INVXLTS
x47INVXLTS n101 w_i1 gnd vdd INVXLTS
x48INVXLTS n103 w_i6 gnd vdd INVXLTS
x49INVXLTS n105 w_i0 gnd vdd INVXLTS
x50INVXLTS n107 w_i7 gnd vdd INVXLTS
x51INVXLTS n109 ld_r gnd vdd INVXLTS
.ends
