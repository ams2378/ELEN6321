
module aes_cipher_top ( clk, rst, ld, done, key, text_in, text_out );
  input [127:0] key;
  input [127:0] text_in;
  output [127:0] text_out;
  input clk, rst, ld;
  output done;
  wire   N21, N32, N33, N34, N35, N36, N37, N38, N39, N48, N49, N50, N51, N52,
         N53, N54, N55, N64, N65, N66, N67, N68, N69, N70, N71, N80, N81, N82,
         N83, N84, N85, N86, N87, N96, N97, N98, N99, N100, N101, N102, N103,
         N112, N113, N114, N115, N116, N117, N118, N119, N128, N129, N130,
         N131, N132, N133, N134, N135, N144, N145, N146, N147, N148, N149,
         N150, N151, N160, N161, N162, N163, N164, N165, N166, N167, N176,
         N177, N178, N179, N180, N181, N182, N183, N192, N193, N194, N195,
         N196, N197, N198, N199, N208, N209, N210, N211, N212, N213, N214,
         N215, N224, N225, N226, N227, N228, N229, N230, N231, N240, N241,
         N242, N243, N244, N245, N246, N247, N256, N257, N258, N259, N260,
         N261, N262, N263, N272, N273, N274, N275, N276, N277, N278, N279,
         N376, N377, N378, N379, N380, N381, N382, N383, N384, N385, N386,
         N387, N388, N389, N390, N391, N392, N393, N394, N395, N396, N397,
         N398, N399, N400, N401, N402, N403, N404, N405, N406, N407, N408,
         N409, N410, N411, N412, N413, N414, N415, N416, N417, N418, N419,
         N420, N421, N422, N423, N424, N425, N426, N427, N428, N429, N430,
         N431, N432, N433, N434, N435, N436, N437, N438, N439, N440, N441,
         N442, N443, N444, N445, N446, N447, N448, N449, N450, N451, N452,
         N453, N454, N455, N456, N457, N458, N459, N460, N461, N462, N463,
         N464, N465, N466, N467, N468, N469, N470, N471, N472, N473, N474,
         N475, N476, N477, N478, N479, N480, N481, N482, N483, N484, N485,
         N486, N487, N488, N489, N490, N491, N492, N493, N494, N495, N496,
         N497, N498, N499, N500, N501, N502, N503, n133, n139, n985, n986,
         n987, n988, n1198, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1266, n1268, n1269, n1270, n1271, n1272, n1273, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1296, n1297, n1298,
         n1299, n1300, n1301, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1327, n1328, n1329, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1447, n1448, n1449, n1450,
         n1451, n1452, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1498, n1499, n1500, n1501, n1502, n1503,
         n1506, n1507, n1508, n1509, n1511, n1512, n1513, n1515, n1516, n1517,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1528, n1529,
         n1531, n1533, n1534, n1535, n1536, n1538, n1540, n1542, n1543, n1544,
         n1546, n1548, n1549, n1550, n1551, n1553, n1555, n1557, n1558, n1560,
         n1562, n1563, n1565, n1566, n1567, n1568, n1569, n1570, n1573, n1574,
         n1576, n1577, n1579, n1580, n1581, n1582, n1583, n1584, n1587, n1588,
         n1590, n1591, n1593, n1594, n1595, n1596, n1597, n1598, n1600, n1601,
         n1602, n1604, n1605, n1607, n1608, n1611, n1612, n1614, n1615, n1616,
         n1618, n1619, n1621, n1622, n1623, n1625, n1626, n1628, n1629, n1630,
         n1632, n1633, n1635, n1637, n1641, n1643, n1644, n1645, n1647, n1648,
         n1650, n1651, n1652, n1653, n1654, n1655, n1659, n1662, n1663, n1665,
         n1667, n1668, n1669, n1670, n1671, n1672, n1674, n1675, n1676, n1682,
         n1683, n1684, n1686, n1687, n1689, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1716, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1773,
         n1774, n1776, n1777, n1778, n1780, n1781, n1783, n1784, n1785, n1787,
         n1788, n1789, n1790, n1791, n1792, n1795, n1796, n1799, n1802, n1803,
         n1804, n1805, n1806, n1807, n1809, n1810, n1811, n1813, n1817, n1819,
         n1820, n1821, n1822, n1823, n1824, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1901, n1902, n1903, n1904, n1905,
         n1906, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1966, n1967, n1968, n1969, n1971, n1972,
         n1974, n1975, n1976, n1977, n1978, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1989, n1991, n1992, n1993, n1995, n1996, n1997,
         n1999, n2000, n2001, n2002, n2006, n2008, n2010, n2012, n2013, n2014,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2029,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2047, n2048, n2053, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2063, n2065, n2066, n2069, n2070, n2073,
         n2074, n2075, n2076, n2079, n2080, n2081, n2083, n2086, n2087, n2088,
         n2089, n2093, n2094, n2095, n2096, n2097, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2149, n2150, n2151, n2152, n2153, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2163, n2164, n2165, n2167, n2168,
         n2169, n2171, n2173, n2178, n2181, n2182, n2185, n2186, n2187, n2188,
         n2189, n2194, n2195, n2196, n2197, n2198, n2199, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2224,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2315, n2316, n2317, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2508, n2509, n2510, n2511, n2512, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2644, n2645, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2835, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2911, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3303, n3305, n3306, n3313, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3488, n3489, n3490, n3492,
         n3493, n3494, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3552, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3618, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3654,
         n3655, n3656, n3657, n3659, n3660, n3661, n3662, n3663, n3665, n3666,
         n3667, n3668, n3671, n3672, n3673, n3674, n3675, n3681, n3685, n3686,
         n3687, n3688, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3698,
         n3699, n3701, n3702, n3706, n3707, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3747, n3752, n3753, n3754,
         n3756, n3757, n3758, n3760, n3761, n3762, n3764, n3765, n3768, n3772,
         n3773, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3791, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3816, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3835,
         n3837, n3838, n3839, n3841, n3842, n3844, n3846, n3852, n3853, n3854,
         n3856, n3859, n3861, n3862, n3863, n3864, n3865, n3866, n3868, n3869,
         n3870, n3871, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3924, n3925, n3926, n3927, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3937, n3938, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3956, n3960, n3961,
         n3962, n3963, n3966, n3967, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4061, n4062, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4153, n4154, n4155, n4156,
         n4157, n4158, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4477,
         n4478, n4479, n4480, n4481, n4482, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4570, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4635, n4642,
         n4643, n4644, n4645, n4646, n4647, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4738, n4739,
         n4740, n4741, n4742, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4818, n4819, n4822, n4824, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4837, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4856, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4932, n4934,
         n4935, n4936, n4937, n4938, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n5006, n5007, n5008, n5009, n5010, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5286, n5287, n5290, n5291, n5292,
         n5293, n5294, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5457, n5461, n5462, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5523, n5527, n5528, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5546,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5611, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5630, n5632, n5633, n5634, n5637, n5639, n5641, n5643, n5644,
         n5648, n5650, n5652, n5655, n5657, n5658, n5660, n5661, n5662, n5663,
         n5664, n5668, n5669, n5670, n5671, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5861, n5862, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5917, n5918, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5968, n5969, n5970, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5997, n5998, n5999, n6000, n6001, n6002, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6063, n6064, n6065, n6066, n6067,
         n6068, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6107, n6108, n6109, n6110,
         n6111, n6112, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6507, n6514, n6515, n6516, n6517,
         n6518, n6519, n6521, n6522, n6531, n6532, n6533, n6534, n6542, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6616,
         n6617, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6655, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6691, n6692, n6693,
         n6694, n6695, n6696, n6699, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6731, n6733, n6734, n6735, n6736, n6737, n6738,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6805, n6806, n6807,
         n6808, n6809, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7130, n7131, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7182, n7183,
         n7184, n7185, n7186, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7240, n7241, n7242, n7243, n7244, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7255, n7256, n7259, n7261, n7262, n7263, n7264,
         n7265, n7268, n7269, n7270, n7273, n7275, n7276, n7280, n7281, n7285,
         n7286, n7289, n7291, n7292, n7293, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7378, n7379, n7380, n7381, n7382, n7383,
         n7385, n7386, n7387, n7388, n7389, n7390, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7406,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7491, n7492,
         n7493, n7494, n7495, n7496, n7498, n7499, n7500, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7528, n7529, n7530, n7531, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7556, n7560, n7561, n7562, n7563, n7564,
         n7567, n7568, n7569, n7570, n7574, n7575, n7576, n7578, n7582, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7607, n7608, n7610, n7611, n7612, n7613, n7615, n7616, n7617, n7618,
         n7619, n7621, n7622, n7625, n7627, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7677, n7679, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7746, n7753, n7754, n7755, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7860, n7861,
         n7865, n7870, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8175, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8261, n8262, n8263, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8291, n8292, n8293, n8294, n8295, n8296, n8301, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8351, n8352,
         n8353, n8354, n8358, n8362, n8363, n8364, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8607,
         n8608, n8609, n8610, n8611, n8612, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8672, n8673, n8674, n8675, n8676, n8677, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765;
  wire   [3:0] dcnt;
  wire   [127:0] text_in_r;
  wire   [31:0] w3;
  wire   [7:0] sa33;
  wire   [7:0] sa23;
  wire   [7:0] sa13;
  wire   [7:0] sa03;
  wire   [31:0] w2;
  wire   [7:0] sa32;
  wire   [7:0] sa22;
  wire   [7:0] sa12;
  wire   [7:0] sa02;
  wire   [31:0] w1;
  wire   [7:0] sa31;
  wire   [7:0] sa21;
  wire   [7:0] sa11;
  wire   [7:0] sa01;
  wire   [31:0] w0;
  wire   [7:0] sa30;
  wire   [7:0] sa20;
  wire   [7:0] sa10;
  wire   [7:0] sa00;
  assign n1198 = ld;

  aes_key_expand_128 u0 ( .clk(clk), .kld(n1198), .key(key), .wo_0(w0), .wo_1(
        w1), .wo_2(w2), .wo_3(w3) );
  EDFFX1TS \text_in_r_reg[127]  ( .D(text_in[127]), .E(n11659), .CK(clk), .Q(
        text_in_r[127]) );
  EDFFX1TS \text_in_r_reg[126]  ( .D(text_in[126]), .E(n11961), .CK(clk), .Q(
        text_in_r[126]) );
  EDFFX1TS \text_in_r_reg[125]  ( .D(text_in[125]), .E(n11657), .CK(clk), .Q(
        text_in_r[125]) );
  EDFFX1TS \text_in_r_reg[124]  ( .D(text_in[124]), .E(n10365), .CK(clk), .Q(
        text_in_r[124]) );
  EDFFX1TS \text_in_r_reg[123]  ( .D(text_in[123]), .E(n11968), .CK(clk), .Q(
        text_in_r[123]) );
  EDFFX1TS \text_in_r_reg[122]  ( .D(text_in[122]), .E(n11658), .CK(clk), .Q(
        text_in_r[122]) );
  EDFFX1TS \text_in_r_reg[121]  ( .D(text_in[121]), .E(n11657), .CK(clk), .Q(
        text_in_r[121]) );
  EDFFX1TS \text_in_r_reg[120]  ( .D(text_in[120]), .E(n10365), .CK(clk), .Q(
        text_in_r[120]) );
  EDFFX1TS \text_in_r_reg[119]  ( .D(text_in[119]), .E(n10361), .CK(clk), .Q(
        text_in_r[119]) );
  EDFFX1TS \text_in_r_reg[118]  ( .D(text_in[118]), .E(n9041), .CK(clk), .Q(
        text_in_r[118]) );
  EDFFX1TS \text_in_r_reg[117]  ( .D(text_in[117]), .E(n11964), .CK(clk), .Q(
        text_in_r[117]) );
  EDFFX1TS \text_in_r_reg[116]  ( .D(text_in[116]), .E(n11664), .CK(clk), .Q(
        text_in_r[116]) );
  EDFFX1TS \text_in_r_reg[115]  ( .D(text_in[115]), .E(n11650), .CK(clk), .Q(
        text_in_r[115]) );
  EDFFX1TS \text_in_r_reg[114]  ( .D(text_in[114]), .E(n12655), .CK(clk), .Q(
        text_in_r[114]) );
  EDFFX1TS \text_in_r_reg[113]  ( .D(text_in[113]), .E(n11657), .CK(clk), .Q(
        text_in_r[113]) );
  EDFFX1TS \text_in_r_reg[112]  ( .D(text_in[112]), .E(n10362), .CK(clk), .Q(
        text_in_r[112]) );
  EDFFX1TS \text_in_r_reg[111]  ( .D(text_in[111]), .E(n11657), .CK(clk), .Q(
        text_in_r[111]) );
  EDFFX1TS \text_in_r_reg[110]  ( .D(text_in[110]), .E(n10366), .CK(clk), .Q(
        text_in_r[110]) );
  EDFFX1TS \text_in_r_reg[109]  ( .D(text_in[109]), .E(n11649), .CK(clk), .Q(
        text_in_r[109]) );
  EDFFX1TS \text_in_r_reg[108]  ( .D(text_in[108]), .E(n10362), .CK(clk), .Q(
        text_in_r[108]) );
  EDFFX1TS \text_in_r_reg[107]  ( .D(text_in[107]), .E(n12607), .CK(clk), .Q(
        text_in_r[107]) );
  EDFFX1TS \text_in_r_reg[106]  ( .D(text_in[106]), .E(n11649), .CK(clk), .Q(
        text_in_r[106]) );
  EDFFX1TS \text_in_r_reg[105]  ( .D(text_in[105]), .E(n12608), .CK(clk), .Q(
        text_in_r[105]) );
  EDFFX1TS \text_in_r_reg[104]  ( .D(text_in[104]), .E(n12606), .CK(clk), .Q(
        text_in_r[104]) );
  EDFFX1TS \text_in_r_reg[103]  ( .D(text_in[103]), .E(n11651), .CK(clk), .Q(
        text_in_r[103]) );
  EDFFX1TS \text_in_r_reg[102]  ( .D(text_in[102]), .E(n11651), .CK(clk), .Q(
        text_in_r[102]) );
  EDFFX1TS \text_in_r_reg[101]  ( .D(text_in[101]), .E(n11965), .CK(clk), .Q(
        text_in_r[101]) );
  EDFFX1TS \text_in_r_reg[100]  ( .D(text_in[100]), .E(n12608), .CK(clk), .Q(
        text_in_r[100]) );
  EDFFX1TS \text_in_r_reg[99]  ( .D(text_in[99]), .E(n11663), .CK(clk), .Q(
        text_in_r[99]) );
  EDFFX1TS \text_in_r_reg[98]  ( .D(text_in[98]), .E(n10362), .CK(clk), .Q(
        text_in_r[98]) );
  EDFFX1TS \text_in_r_reg[97]  ( .D(text_in[97]), .E(n11963), .CK(clk), .Q(
        text_in_r[97]) );
  EDFFX1TS \text_in_r_reg[96]  ( .D(text_in[96]), .E(n11649), .CK(clk), .Q(
        text_in_r[96]) );
  EDFFX1TS \text_in_r_reg[95]  ( .D(text_in[95]), .E(n9041), .CK(clk), .Q(
        text_in_r[95]) );
  EDFFX1TS \text_in_r_reg[94]  ( .D(text_in[94]), .E(n11656), .CK(clk), .Q(
        text_in_r[94]) );
  EDFFX1TS \text_in_r_reg[93]  ( .D(text_in[93]), .E(n11963), .CK(clk), .Q(
        text_in_r[93]) );
  EDFFX1TS \text_in_r_reg[92]  ( .D(text_in[92]), .E(n11656), .CK(clk), .Q(
        text_in_r[92]) );
  EDFFX1TS \text_in_r_reg[91]  ( .D(text_in[91]), .E(n11651), .CK(clk), .Q(
        text_in_r[91]) );
  EDFFX1TS \text_in_r_reg[90]  ( .D(text_in[90]), .E(n9041), .CK(clk), .Q(
        text_in_r[90]) );
  EDFFX1TS \text_in_r_reg[89]  ( .D(text_in[89]), .E(n11665), .CK(clk), .Q(
        text_in_r[89]) );
  EDFFX1TS \text_in_r_reg[88]  ( .D(text_in[88]), .E(n11965), .CK(clk), .Q(
        text_in_r[88]) );
  EDFFX1TS \text_in_r_reg[87]  ( .D(text_in[87]), .E(n11964), .CK(clk), .Q(
        text_in_r[87]) );
  EDFFX1TS \text_in_r_reg[86]  ( .D(text_in[86]), .E(n11961), .CK(clk), .Q(
        text_in_r[86]) );
  EDFFX1TS \text_in_r_reg[85]  ( .D(text_in[85]), .E(n11969), .CK(clk), .Q(
        text_in_r[85]) );
  EDFFX1TS \text_in_r_reg[84]  ( .D(text_in[84]), .E(n12609), .CK(clk), .Q(
        text_in_r[84]) );
  EDFFX1TS \text_in_r_reg[83]  ( .D(text_in[83]), .E(n10365), .CK(clk), .Q(
        text_in_r[83]) );
  EDFFX1TS \text_in_r_reg[82]  ( .D(text_in[82]), .E(n11968), .CK(clk), .Q(
        text_in_r[82]) );
  EDFFX1TS \text_in_r_reg[81]  ( .D(text_in[81]), .E(n12608), .CK(clk), .Q(
        text_in_r[81]) );
  EDFFX1TS \text_in_r_reg[80]  ( .D(text_in[80]), .E(n12609), .CK(clk), .Q(
        text_in_r[80]) );
  EDFFX1TS \text_in_r_reg[79]  ( .D(text_in[79]), .E(n11665), .CK(clk), .Q(
        text_in_r[79]) );
  EDFFX1TS \text_in_r_reg[78]  ( .D(text_in[78]), .E(n11665), .CK(clk), .Q(
        text_in_r[78]) );
  EDFFX1TS \text_in_r_reg[77]  ( .D(text_in[77]), .E(n11666), .CK(clk), .Q(
        text_in_r[77]) );
  EDFFX1TS \text_in_r_reg[76]  ( .D(text_in[76]), .E(n11961), .CK(clk), .Q(
        text_in_r[76]) );
  EDFFX1TS \text_in_r_reg[75]  ( .D(text_in[75]), .E(n11968), .CK(clk), .Q(
        text_in_r[75]) );
  EDFFX1TS \text_in_r_reg[74]  ( .D(text_in[74]), .E(n11960), .CK(clk), .Q(
        text_in_r[74]) );
  EDFFX1TS \text_in_r_reg[73]  ( .D(text_in[73]), .E(n11960), .CK(clk), .Q(
        text_in_r[73]) );
  EDFFX1TS \text_in_r_reg[72]  ( .D(text_in[72]), .E(n11962), .CK(clk), .Q(
        text_in_r[72]) );
  EDFFX1TS \text_in_r_reg[71]  ( .D(text_in[71]), .E(n11967), .CK(clk), .Q(
        text_in_r[71]) );
  EDFFX1TS \text_in_r_reg[70]  ( .D(text_in[70]), .E(n10366), .CK(clk), .Q(
        text_in_r[70]) );
  EDFFX1TS \text_in_r_reg[69]  ( .D(text_in[69]), .E(n11967), .CK(clk), .Q(
        text_in_r[69]) );
  EDFFX1TS \text_in_r_reg[68]  ( .D(text_in[68]), .E(n11961), .CK(clk), .Q(
        text_in_r[68]) );
  EDFFX1TS \text_in_r_reg[67]  ( .D(text_in[67]), .E(n11663), .CK(clk), .Q(
        text_in_r[67]) );
  EDFFX1TS \text_in_r_reg[66]  ( .D(text_in[66]), .E(n11661), .CK(clk), .Q(
        text_in_r[66]) );
  EDFFX1TS \text_in_r_reg[65]  ( .D(text_in[65]), .E(n11661), .CK(clk), .Q(
        text_in_r[65]) );
  EDFFX1TS \text_in_r_reg[64]  ( .D(text_in[64]), .E(n11969), .CK(clk), .Q(
        text_in_r[64]) );
  EDFFX1TS \text_in_r_reg[63]  ( .D(text_in[63]), .E(n12609), .CK(clk), .Q(
        text_in_r[63]) );
  EDFFX1TS \text_in_r_reg[62]  ( .D(text_in[62]), .E(n11960), .CK(clk), .Q(
        text_in_r[62]) );
  EDFFX1TS \text_in_r_reg[61]  ( .D(text_in[61]), .E(n11960), .CK(clk), .Q(
        text_in_r[61]) );
  EDFFX1TS \text_in_r_reg[60]  ( .D(text_in[60]), .E(n11659), .CK(clk), .Q(
        text_in_r[60]) );
  EDFFX1TS \text_in_r_reg[59]  ( .D(text_in[59]), .E(n11659), .CK(clk), .Q(
        text_in_r[59]) );
  EDFFX1TS \text_in_r_reg[58]  ( .D(text_in[58]), .E(n12610), .CK(clk), .Q(
        text_in_r[58]) );
  EDFFX1TS \text_in_r_reg[57]  ( .D(text_in[57]), .E(n11965), .CK(clk), .Q(
        text_in_r[57]) );
  EDFFX1TS \text_in_r_reg[56]  ( .D(text_in[56]), .E(n11660), .CK(clk), .Q(
        text_in_r[56]) );
  EDFFX1TS \text_in_r_reg[55]  ( .D(text_in[55]), .E(n11660), .CK(clk), .Q(
        text_in_r[55]) );
  EDFFX1TS \text_in_r_reg[54]  ( .D(text_in[54]), .E(n11661), .CK(clk), .Q(
        text_in_r[54]) );
  EDFFX1TS \text_in_r_reg[53]  ( .D(text_in[53]), .E(n11660), .CK(clk), .Q(
        text_in_r[53]) );
  EDFFX1TS \text_in_r_reg[52]  ( .D(text_in[52]), .E(n11963), .CK(clk), .Q(
        text_in_r[52]) );
  EDFFX1TS \text_in_r_reg[51]  ( .D(text_in[51]), .E(n12609), .CK(clk), .Q(
        text_in_r[51]) );
  EDFFX1TS \text_in_r_reg[50]  ( .D(text_in[50]), .E(n11963), .CK(clk), .Q(
        text_in_r[50]) );
  EDFFX1TS \text_in_r_reg[49]  ( .D(text_in[49]), .E(n11663), .CK(clk), .Q(
        text_in_r[49]) );
  EDFFX1TS \text_in_r_reg[48]  ( .D(text_in[48]), .E(n12607), .CK(clk), .Q(
        text_in_r[48]) );
  EDFFX1TS \text_in_r_reg[47]  ( .D(text_in[47]), .E(n11962), .CK(clk), .Q(
        text_in_r[47]) );
  EDFFX1TS \text_in_r_reg[46]  ( .D(text_in[46]), .E(n11969), .CK(clk), .Q(
        text_in_r[46]) );
  EDFFX1TS \text_in_r_reg[45]  ( .D(text_in[45]), .E(n11967), .CK(clk), .Q(
        text_in_r[45]) );
  EDFFX1TS \text_in_r_reg[44]  ( .D(text_in[44]), .E(n11962), .CK(clk), .Q(
        text_in_r[44]) );
  EDFFX1TS \text_in_r_reg[43]  ( .D(text_in[43]), .E(n11967), .CK(clk), .Q(
        text_in_r[43]) );
  EDFFX1TS \text_in_r_reg[42]  ( .D(text_in[42]), .E(n11667), .CK(clk), .Q(
        text_in_r[42]) );
  EDFFX1TS \text_in_r_reg[41]  ( .D(text_in[41]), .E(n11962), .CK(clk), .Q(
        text_in_r[41]) );
  EDFFX1TS \text_in_r_reg[40]  ( .D(text_in[40]), .E(n11667), .CK(clk), .Q(
        text_in_r[40]) );
  EDFFX1TS \text_in_r_reg[39]  ( .D(text_in[39]), .E(n11650), .CK(clk), .Q(
        text_in_r[39]) );
  EDFFX1TS \text_in_r_reg[38]  ( .D(text_in[38]), .E(n11964), .CK(clk), .Q(
        text_in_r[38]) );
  EDFFX1TS \text_in_r_reg[37]  ( .D(text_in[37]), .E(n11665), .CK(clk), .Q(
        text_in_r[37]) );
  EDFFX1TS \text_in_r_reg[36]  ( .D(text_in[36]), .E(n11968), .CK(clk), .Q(
        text_in_r[36]) );
  EDFFX1TS \text_in_r_reg[35]  ( .D(text_in[35]), .E(n11667), .CK(clk), .Q(
        text_in_r[35]) );
  EDFFX1TS \text_in_r_reg[34]  ( .D(text_in[34]), .E(n11649), .CK(clk), .Q(
        text_in_r[34]) );
  EDFFX1TS \text_in_r_reg[33]  ( .D(text_in[33]), .E(n10361), .CK(clk), .Q(
        text_in_r[33]) );
  EDFFX1TS \text_in_r_reg[32]  ( .D(text_in[32]), .E(n11666), .CK(clk), .Q(
        text_in_r[32]) );
  EDFFX1TS \text_in_r_reg[31]  ( .D(text_in[31]), .E(n11661), .CK(clk), .Q(
        text_in_r[31]) );
  EDFFX1TS \text_in_r_reg[30]  ( .D(text_in[30]), .E(n11663), .CK(clk), .Q(
        text_in_r[30]) );
  EDFFX1TS \text_in_r_reg[29]  ( .D(text_in[29]), .E(n10366), .CK(clk), .Q(
        text_in_r[29]) );
  EDFFX1TS \text_in_r_reg[28]  ( .D(text_in[28]), .E(n11658), .CK(clk), .Q(
        text_in_r[28]) );
  EDFFX1TS \text_in_r_reg[27]  ( .D(text_in[27]), .E(n11666), .CK(clk), .Q(
        text_in_r[27]) );
  EDFFX1TS \text_in_r_reg[26]  ( .D(text_in[26]), .E(n12610), .CK(clk), .Q(
        text_in_r[26]) );
  EDFFX1TS \text_in_r_reg[25]  ( .D(text_in[25]), .E(n11658), .CK(clk), .Q(
        text_in_r[25]) );
  EDFFX1TS \text_in_r_reg[24]  ( .D(text_in[24]), .E(n11656), .CK(clk), .Q(
        text_in_r[24]) );
  EDFFX1TS \text_in_r_reg[23]  ( .D(text_in[23]), .E(n12610), .CK(clk), .Q(
        text_in_r[23]) );
  EDFFX1TS \text_in_r_reg[22]  ( .D(text_in[22]), .E(n12607), .CK(clk), .Q(
        text_in_r[22]) );
  EDFFX1TS \text_in_r_reg[21]  ( .D(text_in[21]), .E(n10365), .CK(clk), .Q(
        text_in_r[21]) );
  EDFFX1TS \text_in_r_reg[20]  ( .D(text_in[20]), .E(n11667), .CK(clk), .Q(
        text_in_r[20]) );
  EDFFX1TS \text_in_r_reg[19]  ( .D(text_in[19]), .E(n11656), .CK(clk), .Q(
        text_in_r[19]) );
  EDFFX1TS \text_in_r_reg[18]  ( .D(text_in[18]), .E(n11964), .CK(clk), .Q(
        text_in_r[18]) );
  EDFFX1TS \text_in_r_reg[17]  ( .D(text_in[17]), .E(n11666), .CK(clk), .Q(
        text_in_r[17]) );
  EDFFX1TS \text_in_r_reg[16]  ( .D(text_in[16]), .E(n11650), .CK(clk), .Q(
        text_in_r[16]) );
  EDFFX1TS \text_in_r_reg[15]  ( .D(text_in[15]), .E(n12610), .CK(clk), .Q(
        text_in_r[15]) );
  EDFFX1TS \text_in_r_reg[14]  ( .D(text_in[14]), .E(n11664), .CK(clk), .Q(
        text_in_r[14]) );
  EDFFX1TS \text_in_r_reg[13]  ( .D(text_in[13]), .E(n10361), .CK(clk), .Q(
        text_in_r[13]) );
  EDFFX1TS \text_in_r_reg[12]  ( .D(text_in[12]), .E(n11658), .CK(clk), .Q(
        text_in_r[12]) );
  EDFFX1TS \text_in_r_reg[11]  ( .D(text_in[11]), .E(n12611), .CK(clk), .Q(
        text_in_r[11]) );
  EDFFX1TS \text_in_r_reg[10]  ( .D(text_in[10]), .E(n10362), .CK(clk), .Q(
        text_in_r[10]) );
  EDFFX1TS \text_in_r_reg[9]  ( .D(text_in[9]), .E(n10361), .CK(clk), .Q(
        text_in_r[9]) );
  EDFFX1TS \text_in_r_reg[8]  ( .D(text_in[8]), .E(n11651), .CK(clk), .Q(
        text_in_r[8]) );
  EDFFX1TS \text_in_r_reg[7]  ( .D(text_in[7]), .E(n12612), .CK(clk), .Q(
        text_in_r[7]) );
  EDFFX1TS \text_in_r_reg[6]  ( .D(text_in[6]), .E(n11664), .CK(clk), .Q(
        text_in_r[6]) );
  EDFFX1TS \text_in_r_reg[5]  ( .D(text_in[5]), .E(n11650), .CK(clk), .Q(
        text_in_r[5]) );
  EDFFX1TS \text_in_r_reg[4]  ( .D(text_in[4]), .E(n12606), .CK(clk), .Q(
        text_in_r[4]) );
  EDFFX1TS \text_in_r_reg[3]  ( .D(text_in[3]), .E(n12611), .CK(clk), .Q(
        text_in_r[3]) );
  EDFFX1TS \text_in_r_reg[2]  ( .D(text_in[2]), .E(n11664), .CK(clk), .Q(
        text_in_r[2]) );
  EDFFX1TS \text_in_r_reg[1]  ( .D(text_in[1]), .E(n11660), .CK(clk), .Q(
        text_in_r[1]) );
  EDFFX1TS \text_in_r_reg[0]  ( .D(text_in[0]), .E(n11659), .CK(clk), .Q(
        text_in_r[0]) );
  DFFXLTS \dcnt_reg[3]  ( .D(n987), .CK(clk), .QN(n139) );
  DFFQX1TS done_reg ( .D(N21), .CK(clk), .Q(done) );
  DFFQX1TS \dcnt_reg[1]  ( .D(n986), .CK(clk), .Q(dcnt[1]) );
  DFFQX1TS \text_out_reg[96]  ( .D(N479), .CK(clk), .Q(text_out[96]) );
  DFFQX1TS \text_out_reg[64]  ( .D(N487), .CK(clk), .Q(text_out[64]) );
  DFFQX1TS \text_out_reg[40]  ( .D(N463), .CK(clk), .Q(text_out[40]) );
  DFFQX1TS \text_out_reg[0]  ( .D(N503), .CK(clk), .Q(text_out[0]) );
  DFFQX1TS \text_out_reg[26]  ( .D(N405), .CK(clk), .Q(text_out[26]) );
  DFFQX1TS \text_out_reg[112]  ( .D(N415), .CK(clk), .Q(text_out[112]) );
  DFFQX1TS \text_out_reg[80]  ( .D(N423), .CK(clk), .Q(text_out[80]) );
  DFFQX1TS \text_out_reg[32]  ( .D(N495), .CK(clk), .Q(text_out[32]) );
  DFFQX1TS \text_out_reg[16]  ( .D(N439), .CK(clk), .Q(text_out[16]) );
  DFFQX1TS \text_out_reg[8]  ( .D(N471), .CK(clk), .Q(text_out[8]) );
  DFFQX1TS \text_out_reg[104]  ( .D(N447), .CK(clk), .Q(text_out[104]) );
  DFFQX1TS \text_out_reg[72]  ( .D(N455), .CK(clk), .Q(text_out[72]) );
  DFFQX1TS \text_out_reg[48]  ( .D(N431), .CK(clk), .Q(text_out[48]) );
  DFFQX1TS \text_out_reg[120]  ( .D(N383), .CK(clk), .Q(text_out[120]) );
  DFFQX1TS \text_out_reg[88]  ( .D(N391), .CK(clk), .Q(text_out[88]) );
  DFFQX1TS \text_out_reg[24]  ( .D(N407), .CK(clk), .Q(text_out[24]) );
  DFFQX1TS \text_out_reg[56]  ( .D(N399), .CK(clk), .Q(text_out[56]) );
  DFFQX1TS \text_out_reg[2]  ( .D(N501), .CK(clk), .Q(text_out[2]) );
  DFFQX1TS \text_out_reg[98]  ( .D(N477), .CK(clk), .Q(text_out[98]) );
  DFFQX1TS \text_out_reg[66]  ( .D(N485), .CK(clk), .Q(text_out[66]) );
  DFFQX1TS \text_out_reg[42]  ( .D(N461), .CK(clk), .Q(text_out[42]) );
  DFFQX1TS \text_out_reg[99]  ( .D(N476), .CK(clk), .Q(text_out[99]) );
  DFFQX1TS \text_out_reg[67]  ( .D(N484), .CK(clk), .Q(text_out[67]) );
  DFFQX1TS \text_out_reg[43]  ( .D(N460), .CK(clk), .Q(text_out[43]) );
  DFFQX1TS \text_out_reg[3]  ( .D(N500), .CK(clk), .Q(text_out[3]) );
  DFFQX1TS \text_out_reg[51]  ( .D(N428), .CK(clk), .Q(text_out[51]) );
  DFFQX1TS \text_out_reg[123]  ( .D(N380), .CK(clk), .Q(text_out[123]) );
  DFFQX1TS \text_out_reg[91]  ( .D(N388), .CK(clk), .Q(text_out[91]) );
  DFFQX1TS \text_out_reg[115]  ( .D(N412), .CK(clk), .Q(text_out[115]) );
  DFFQX1TS \text_out_reg[83]  ( .D(N420), .CK(clk), .Q(text_out[83]) );
  DFFQX1TS \text_out_reg[35]  ( .D(N492), .CK(clk), .Q(text_out[35]) );
  DFFQX1TS \text_out_reg[27]  ( .D(N404), .CK(clk), .Q(text_out[27]) );
  DFFQX1TS \text_out_reg[11]  ( .D(N468), .CK(clk), .Q(text_out[11]) );
  DFFQX1TS \text_out_reg[107]  ( .D(N444), .CK(clk), .Q(text_out[107]) );
  DFFQX1TS \text_out_reg[75]  ( .D(N452), .CK(clk), .Q(text_out[75]) );
  DFFQX1TS \text_out_reg[59]  ( .D(N396), .CK(clk), .Q(text_out[59]) );
  DFFQX1TS \text_out_reg[19]  ( .D(N436), .CK(clk), .Q(text_out[19]) );
  DFFQX1TS \text_out_reg[50]  ( .D(N429), .CK(clk), .Q(text_out[50]) );
  DFFQX1TS \text_out_reg[18]  ( .D(N437), .CK(clk), .Q(text_out[18]) );
  DFFQX1TS \text_out_reg[114]  ( .D(N413), .CK(clk), .Q(text_out[114]) );
  DFFQX1TS \text_out_reg[82]  ( .D(N421), .CK(clk), .Q(text_out[82]) );
  DFFQX1TS \text_out_reg[58]  ( .D(N397), .CK(clk), .Q(text_out[58]) );
  DFFQX1TS \text_out_reg[34]  ( .D(N493), .CK(clk), .Q(text_out[34]) );
  DFFQX1TS \text_out_reg[10]  ( .D(N469), .CK(clk), .Q(text_out[10]) );
  DFFQX1TS \text_out_reg[106]  ( .D(N445), .CK(clk), .Q(text_out[106]) );
  DFFQX1TS \text_out_reg[74]  ( .D(N453), .CK(clk), .Q(text_out[74]) );
  DFFQX1TS \text_out_reg[122]  ( .D(N381), .CK(clk), .Q(text_out[122]) );
  DFFQX1TS \text_out_reg[90]  ( .D(N389), .CK(clk), .Q(text_out[90]) );
  DFFQX1TS \text_out_reg[30]  ( .D(N401), .CK(clk), .Q(text_out[30]) );
  DFFQX1TS \text_out_reg[29]  ( .D(N402), .CK(clk), .Q(text_out[29]) );
  DFFQX1TS \text_out_reg[6]  ( .D(N497), .CK(clk), .Q(text_out[6]) );
  DFFQX1TS \text_out_reg[102]  ( .D(N473), .CK(clk), .Q(text_out[102]) );
  DFFQX1TS \text_out_reg[70]  ( .D(N481), .CK(clk), .Q(text_out[70]) );
  DFFQX1TS \text_out_reg[38]  ( .D(N489), .CK(clk), .Q(text_out[38]) );
  DFFQX1TS \text_out_reg[41]  ( .D(N462), .CK(clk), .Q(text_out[41]) );
  DFFQX1TS \text_out_reg[125]  ( .D(N378), .CK(clk), .Q(text_out[125]) );
  DFFQX1TS \text_out_reg[93]  ( .D(N386), .CK(clk), .Q(text_out[93]) );
  DFFQX1TS \text_out_reg[61]  ( .D(N394), .CK(clk), .Q(text_out[61]) );
  DFFQX1TS \text_out_reg[5]  ( .D(N498), .CK(clk), .Q(text_out[5]) );
  DFFQX1TS \text_out_reg[100]  ( .D(N475), .CK(clk), .Q(text_out[100]) );
  DFFQX1TS \text_out_reg[68]  ( .D(N483), .CK(clk), .Q(text_out[68]) );
  DFFQX1TS \text_out_reg[118]  ( .D(N409), .CK(clk), .Q(text_out[118]) );
  DFFQX1TS \text_out_reg[86]  ( .D(N417), .CK(clk), .Q(text_out[86]) );
  DFFQX1TS \text_out_reg[54]  ( .D(N425), .CK(clk), .Q(text_out[54]) );
  DFFQX1TS \text_out_reg[14]  ( .D(N465), .CK(clk), .Q(text_out[14]) );
  DFFQX1TS \text_out_reg[36]  ( .D(N491), .CK(clk), .Q(text_out[36]) );
  DFFQX1TS \text_out_reg[4]  ( .D(N499), .CK(clk), .Q(text_out[4]) );
  DFFQX1TS \text_out_reg[110]  ( .D(N441), .CK(clk), .Q(text_out[110]) );
  DFFQX1TS \text_out_reg[78]  ( .D(N449), .CK(clk), .Q(text_out[78]) );
  DFFQX1TS \text_out_reg[46]  ( .D(N457), .CK(clk), .Q(text_out[46]) );
  DFFQX1TS \text_out_reg[22]  ( .D(N433), .CK(clk), .Q(text_out[22]) );
  DFFQX1TS \text_out_reg[126]  ( .D(N377), .CK(clk), .Q(text_out[126]) );
  DFFQX1TS \text_out_reg[94]  ( .D(N385), .CK(clk), .Q(text_out[94]) );
  DFFQX1TS \text_out_reg[62]  ( .D(N393), .CK(clk), .Q(text_out[62]) );
  DFFQX1TS \text_out_reg[97]  ( .D(N478), .CK(clk), .Q(text_out[97]) );
  DFFQX1TS \text_out_reg[65]  ( .D(N486), .CK(clk), .Q(text_out[65]) );
  DFFQX1TS \text_out_reg[1]  ( .D(N502), .CK(clk), .Q(text_out[1]) );
  DFFQX1TS \text_out_reg[101]  ( .D(N474), .CK(clk), .Q(text_out[101]) );
  DFFQX1TS \text_out_reg[69]  ( .D(N482), .CK(clk), .Q(text_out[69]) );
  DFFQX1TS \text_out_reg[37]  ( .D(N490), .CK(clk), .Q(text_out[37]) );
  DFFQX1TS \text_out_reg[124]  ( .D(N379), .CK(clk), .Q(text_out[124]) );
  DFFQX1TS \text_out_reg[92]  ( .D(N387), .CK(clk), .Q(text_out[92]) );
  DFFQX1TS \text_out_reg[60]  ( .D(N395), .CK(clk), .Q(text_out[60]) );
  DFFQX1TS \text_out_reg[121]  ( .D(N382), .CK(clk), .Q(text_out[121]) );
  DFFQX1TS \text_out_reg[89]  ( .D(N390), .CK(clk), .Q(text_out[89]) );
  DFFQX1TS \text_out_reg[116]  ( .D(N411), .CK(clk), .Q(text_out[116]) );
  DFFQX1TS \text_out_reg[84]  ( .D(N419), .CK(clk), .Q(text_out[84]) );
  DFFQX1TS \text_out_reg[52]  ( .D(N427), .CK(clk), .Q(text_out[52]) );
  DFFQX1TS \text_out_reg[20]  ( .D(N435), .CK(clk), .Q(text_out[20]) );
  DFFQX1TS \text_out_reg[12]  ( .D(N467), .CK(clk), .Q(text_out[12]) );
  DFFQX1TS \text_out_reg[108]  ( .D(N443), .CK(clk), .Q(text_out[108]) );
  DFFQX1TS \text_out_reg[76]  ( .D(N451), .CK(clk), .Q(text_out[76]) );
  DFFQX1TS \text_out_reg[44]  ( .D(N459), .CK(clk), .Q(text_out[44]) );
  DFFQX1TS \text_out_reg[28]  ( .D(N403), .CK(clk), .Q(text_out[28]) );
  DFFQX1TS \text_out_reg[113]  ( .D(N414), .CK(clk), .Q(text_out[113]) );
  DFFQX1TS \text_out_reg[81]  ( .D(N422), .CK(clk), .Q(text_out[81]) );
  DFFQX1TS \text_out_reg[57]  ( .D(N398), .CK(clk), .Q(text_out[57]) );
  DFFQX1TS \text_out_reg[49]  ( .D(N430), .CK(clk), .Q(text_out[49]) );
  DFFQX1TS \text_out_reg[33]  ( .D(N494), .CK(clk), .Q(text_out[33]) );
  DFFQX1TS \text_out_reg[9]  ( .D(N470), .CK(clk), .Q(text_out[9]) );
  DFFQX1TS \text_out_reg[105]  ( .D(N446), .CK(clk), .Q(text_out[105]) );
  DFFQX1TS \text_out_reg[73]  ( .D(N454), .CK(clk), .Q(text_out[73]) );
  DFFQX1TS \text_out_reg[25]  ( .D(N406), .CK(clk), .Q(text_out[25]) );
  DFFQX1TS \text_out_reg[17]  ( .D(N438), .CK(clk), .Q(text_out[17]) );
  DFFQX1TS \text_out_reg[117]  ( .D(N410), .CK(clk), .Q(text_out[117]) );
  DFFQX1TS \text_out_reg[85]  ( .D(N418), .CK(clk), .Q(text_out[85]) );
  DFFQX1TS \text_out_reg[53]  ( .D(N426), .CK(clk), .Q(text_out[53]) );
  DFFQX1TS \text_out_reg[21]  ( .D(N434), .CK(clk), .Q(text_out[21]) );
  DFFQX1TS \text_out_reg[13]  ( .D(N466), .CK(clk), .Q(text_out[13]) );
  DFFQX1TS \text_out_reg[109]  ( .D(N442), .CK(clk), .Q(text_out[109]) );
  DFFQX1TS \text_out_reg[77]  ( .D(N450), .CK(clk), .Q(text_out[77]) );
  DFFQX1TS \text_out_reg[45]  ( .D(N458), .CK(clk), .Q(text_out[45]) );
  DFFQX1TS \text_out_reg[31]  ( .D(N400), .CK(clk), .Q(text_out[31]) );
  DFFQX1TS \text_out_reg[119]  ( .D(N408), .CK(clk), .Q(text_out[119]) );
  DFFQX1TS \text_out_reg[87]  ( .D(N416), .CK(clk), .Q(text_out[87]) );
  DFFQX1TS \text_out_reg[55]  ( .D(N424), .CK(clk), .Q(text_out[55]) );
  DFFQX1TS \text_out_reg[23]  ( .D(N432), .CK(clk), .Q(text_out[23]) );
  DFFQX1TS \text_out_reg[127]  ( .D(N376), .CK(clk), .Q(text_out[127]) );
  DFFQX1TS \text_out_reg[111]  ( .D(N440), .CK(clk), .Q(text_out[111]) );
  DFFQX1TS \text_out_reg[95]  ( .D(N384), .CK(clk), .Q(text_out[95]) );
  DFFQX1TS \text_out_reg[79]  ( .D(N448), .CK(clk), .Q(text_out[79]) );
  DFFQX1TS \text_out_reg[63]  ( .D(N392), .CK(clk), .Q(text_out[63]) );
  DFFQX1TS \text_out_reg[47]  ( .D(N456), .CK(clk), .Q(text_out[47]) );
  DFFQX1TS \text_out_reg[15]  ( .D(N464), .CK(clk), .Q(text_out[15]) );
  DFFQX1TS \text_out_reg[103]  ( .D(N472), .CK(clk), .Q(text_out[103]) );
  DFFQX1TS \text_out_reg[71]  ( .D(N480), .CK(clk), .Q(text_out[71]) );
  DFFQX1TS \text_out_reg[39]  ( .D(N488), .CK(clk), .Q(text_out[39]) );
  DFFQX1TS \text_out_reg[7]  ( .D(N496), .CK(clk), .Q(text_out[7]) );
  DFFQX1TS \sa03_reg[2]  ( .D(N82), .CK(clk), .Q(sa03[2]) );
  DFFQX1TS \sa01_reg[2]  ( .D(N210), .CK(clk), .Q(sa01[2]) );
  DFFQX1TS \sa00_reg[2]  ( .D(N274), .CK(clk), .Q(sa00[2]) );
  DFFQX1TS \sa03_reg[6]  ( .D(N86), .CK(clk), .Q(sa03[6]) );
  DFFQX1TS \sa03_reg[5]  ( .D(N85), .CK(clk), .Q(sa03[5]) );
  DFFQX1TS \sa21_reg[2]  ( .D(N178), .CK(clk), .Q(sa21[2]) );
  DFFQX1TS \sa20_reg[2]  ( .D(N242), .CK(clk), .Q(sa20[2]) );
  DFFQX1TS \sa02_reg[2]  ( .D(N146), .CK(clk), .Q(sa02[2]) );
  DFFQX1TS \sa33_reg[0]  ( .D(N32), .CK(clk), .Q(sa33[0]) );
  DFFQX1TS \sa31_reg[0]  ( .D(N160), .CK(clk), .Q(sa31[0]) );
  DFFQX1TS \sa30_reg[0]  ( .D(N224), .CK(clk), .Q(sa30[0]) );
  DFFQX1TS \sa32_reg[3]  ( .D(N99), .CK(clk), .Q(sa32[3]) );
  DFFQX1TS \sa32_reg[1]  ( .D(N97), .CK(clk), .Q(sa32[1]) );
  DFFQX1TS \sa31_reg[2]  ( .D(N162), .CK(clk), .Q(sa31[2]) );
  DFFQX1TS \sa30_reg[2]  ( .D(N226), .CK(clk), .Q(sa30[2]) );
  DFFQX1TS \sa33_reg[2]  ( .D(N34), .CK(clk), .Q(sa33[2]) );
  DFFQX1TS \sa32_reg[2]  ( .D(N98), .CK(clk), .Q(sa32[2]) );
  DFFQX1TS \sa13_reg[2]  ( .D(N66), .CK(clk), .Q(sa13[2]) );
  DFFQX1TS \sa10_reg[2]  ( .D(N258), .CK(clk), .Q(sa10[2]) );
  DFFQX1TS \sa12_reg[4]  ( .D(N132), .CK(clk), .Q(sa12[4]) );
  DFFQX1TS \sa11_reg[4]  ( .D(N196), .CK(clk), .Q(sa11[4]) );
  DFFQX1TS \sa11_reg[1]  ( .D(N193), .CK(clk), .Q(sa11[1]) );
  DFFQX1TS \sa10_reg[1]  ( .D(N257), .CK(clk), .Q(sa10[1]) );
  DFFQX1TS \sa12_reg[3]  ( .D(N131), .CK(clk), .Q(sa12[3]) );
  DFFQX1TS \sa11_reg[3]  ( .D(N195), .CK(clk), .Q(sa11[3]) );
  DFFQX1TS \sa10_reg[3]  ( .D(N259), .CK(clk), .Q(sa10[3]) );
  DFFQX1TS \sa12_reg[1]  ( .D(N129), .CK(clk), .Q(sa12[1]) );
  DFFQX1TS \sa13_reg[4]  ( .D(N68), .CK(clk), .Q(sa13[4]) );
  DFFQX1TS \sa13_reg[1]  ( .D(N65), .CK(clk), .Q(sa13[1]) );
  DFFQX1TS \sa31_reg[3]  ( .D(N163), .CK(clk), .Q(sa31[3]) );
  DFFQX1TS \sa01_reg[6]  ( .D(N214), .CK(clk), .Q(sa01[6]) );
  DFFQX1TS \sa00_reg[6]  ( .D(N278), .CK(clk), .Q(sa00[6]) );
  DFFQX1TS \sa02_reg[5]  ( .D(N149), .CK(clk), .Q(sa02[5]) );
  DFFQX1TS \sa01_reg[5]  ( .D(N213), .CK(clk), .Q(sa01[5]) );
  DFFQX1TS \sa00_reg[5]  ( .D(N277), .CK(clk), .Q(sa00[5]) );
  DFFQX1TS \sa12_reg[0]  ( .D(N128), .CK(clk), .Q(sa12[0]) );
  DFFQX1TS \sa11_reg[0]  ( .D(N192), .CK(clk), .Q(sa11[0]) );
  DFFQX1TS \sa10_reg[0]  ( .D(N256), .CK(clk), .Q(sa10[0]) );
  DFFQX1TS \sa13_reg[0]  ( .D(N64), .CK(clk), .Q(sa13[0]) );
  DFFQX1TS \sa22_reg[5]  ( .D(N117), .CK(clk), .Q(sa22[5]) );
  DFFQX1TS \sa21_reg[5]  ( .D(N181), .CK(clk), .Q(sa21[5]) );
  DFFQX1TS \sa20_reg[5]  ( .D(N245), .CK(clk), .Q(sa20[5]) );
  DFFQX1TS \sa12_reg[5]  ( .D(N133), .CK(clk), .Q(sa12[5]) );
  DFFQX1TS \sa11_reg[5]  ( .D(N197), .CK(clk), .Q(sa11[5]) );
  DFFQX1TS \sa10_reg[5]  ( .D(N261), .CK(clk), .Q(sa10[5]) );
  DFFQX1TS \sa23_reg[4]  ( .D(N52), .CK(clk), .Q(sa23[4]) );
  DFFQX1TS \sa23_reg[1]  ( .D(N49), .CK(clk), .Q(sa23[1]) );
  DFFQX1TS \sa23_reg[3]  ( .D(N51), .CK(clk), .Q(sa23[3]) );
  DFFQX1TS \sa33_reg[5]  ( .D(N37), .CK(clk), .Q(sa33[5]) );
  DFFQX1TS \sa21_reg[1]  ( .D(N177), .CK(clk), .Q(sa21[1]) );
  DFFQX1TS \sa20_reg[4]  ( .D(N244), .CK(clk), .Q(sa20[4]) );
  DFFQX1TS \sa20_reg[1]  ( .D(N241), .CK(clk), .Q(sa20[1]) );
  DFFQX1TS \sa21_reg[3]  ( .D(N179), .CK(clk), .Q(sa21[3]) );
  DFFQX1TS \sa22_reg[4]  ( .D(N116), .CK(clk), .Q(sa22[4]) );
  DFFQX1TS \sa22_reg[3]  ( .D(N115), .CK(clk), .Q(sa22[3]) );
  DFFQX1TS \sa32_reg[6]  ( .D(N102), .CK(clk), .Q(sa32[6]) );
  DFFQX1TS \sa31_reg[6]  ( .D(N166), .CK(clk), .Q(sa31[6]) );
  DFFQX1TS \sa30_reg[6]  ( .D(N230), .CK(clk), .Q(sa30[6]) );
  DFFQX1TS \sa01_reg[4]  ( .D(N212), .CK(clk), .Q(sa01[4]) );
  DFFQX1TS \sa01_reg[3]  ( .D(N211), .CK(clk), .Q(sa01[3]) );
  DFFQX1TS \sa01_reg[1]  ( .D(N209), .CK(clk), .Q(sa01[1]) );
  DFFQX1TS \sa00_reg[4]  ( .D(N276), .CK(clk), .Q(sa00[4]) );
  DFFQX1TS \sa00_reg[3]  ( .D(N275), .CK(clk), .Q(sa00[3]) );
  DFFQX1TS \sa00_reg[1]  ( .D(N273), .CK(clk), .Q(sa00[1]) );
  DFFQX1TS \sa03_reg[4]  ( .D(N84), .CK(clk), .Q(sa03[4]) );
  DFFQX1TS \sa03_reg[3]  ( .D(N83), .CK(clk), .Q(sa03[3]) );
  DFFQX1TS \sa03_reg[1]  ( .D(N81), .CK(clk), .Q(sa03[1]) );
  DFFQX1TS \sa02_reg[4]  ( .D(N148), .CK(clk), .Q(sa02[4]) );
  DFFQX1TS \sa32_reg[5]  ( .D(N101), .CK(clk), .Q(sa32[5]) );
  DFFQX1TS \sa31_reg[5]  ( .D(N165), .CK(clk), .Q(sa31[5]) );
  DFFQX1TS \sa30_reg[5]  ( .D(N229), .CK(clk), .Q(sa30[5]) );
  DFFQX1TS \sa23_reg[6]  ( .D(N54), .CK(clk), .Q(sa23[6]) );
  DFFQX1TS \sa22_reg[6]  ( .D(N118), .CK(clk), .Q(sa22[6]) );
  DFFQX1TS \sa21_reg[6]  ( .D(N182), .CK(clk), .Q(sa21[6]) );
  DFFQX1TS \sa20_reg[6]  ( .D(N246), .CK(clk), .Q(sa20[6]) );
  DFFQX1TS \sa12_reg[6]  ( .D(N134), .CK(clk), .Q(sa12[6]) );
  DFFQX1TS \sa11_reg[6]  ( .D(N198), .CK(clk), .Q(sa11[6]) );
  DFFQX1TS \sa10_reg[6]  ( .D(N262), .CK(clk), .Q(sa10[6]) );
  DFFQX1TS \sa23_reg[5]  ( .D(N53), .CK(clk), .Q(sa23[5]) );
  DFFQX1TS \sa13_reg[5]  ( .D(N69), .CK(clk), .Q(sa13[5]) );
  DFFQX1TS \sa23_reg[0]  ( .D(N48), .CK(clk), .Q(sa23[0]) );
  DFFQX1TS \sa21_reg[0]  ( .D(N176), .CK(clk), .Q(sa21[0]) );
  DFFQX1TS \sa20_reg[0]  ( .D(N240), .CK(clk), .Q(sa20[0]) );
  DFFQX1TS \sa32_reg[0]  ( .D(N96), .CK(clk), .Q(sa32[0]) );
  DFFQX1TS \sa33_reg[4]  ( .D(N36), .CK(clk), .Q(sa33[4]) );
  DFFQX1TS \sa31_reg[4]  ( .D(N164), .CK(clk), .Q(sa31[4]) );
  DFFQX1TS \sa30_reg[4]  ( .D(N228), .CK(clk), .Q(sa30[4]) );
  DFFQX1TS \sa32_reg[4]  ( .D(N100), .CK(clk), .Q(sa32[4]) );
  DFFQX1TS \sa33_reg[1]  ( .D(N33), .CK(clk), .Q(sa33[1]) );
  DFFQX1TS \sa31_reg[1]  ( .D(N161), .CK(clk), .Q(sa31[1]) );
  DFFQX1TS \sa30_reg[1]  ( .D(N225), .CK(clk), .Q(sa30[1]) );
  DFFQX1TS \sa22_reg[1]  ( .D(N113), .CK(clk), .Q(sa22[1]) );
  DFFQX1TS \sa22_reg[0]  ( .D(N112), .CK(clk), .Q(sa22[0]) );
  DFFQX1TS \sa01_reg[0]  ( .D(N208), .CK(clk), .Q(sa01[0]) );
  DFFQX1TS \sa03_reg[0]  ( .D(N80), .CK(clk), .Q(sa03[0]) );
  DFFQX1TS \sa02_reg[0]  ( .D(N144), .CK(clk), .Q(sa02[0]) );
  DFFQX1TS \sa00_reg[7]  ( .D(N279), .CK(clk), .Q(sa00[7]) );
  DFFQX1TS \sa10_reg[7]  ( .D(N263), .CK(clk), .Q(sa10[7]) );
  DFFQX1TS \sa20_reg[7]  ( .D(N247), .CK(clk), .Q(sa20[7]) );
  DFFQX1TS \sa11_reg[7]  ( .D(N199), .CK(clk), .Q(sa11[7]) );
  DFFQX1TS \sa21_reg[7]  ( .D(N183), .CK(clk), .Q(sa21[7]) );
  DFFQX1TS \sa31_reg[7]  ( .D(N167), .CK(clk), .Q(sa31[7]) );
  DFFQX1TS \sa02_reg[7]  ( .D(N151), .CK(clk), .Q(sa02[7]) );
  DFFQX1TS \sa12_reg[7]  ( .D(N135), .CK(clk), .Q(sa12[7]) );
  DFFQX1TS \sa22_reg[7]  ( .D(N119), .CK(clk), .Q(sa22[7]) );
  DFFQX1TS \sa32_reg[7]  ( .D(N103), .CK(clk), .Q(sa32[7]) );
  DFFQX1TS \sa03_reg[7]  ( .D(N87), .CK(clk), .Q(sa03[7]) );
  DFFQX1TS \sa13_reg[7]  ( .D(N71), .CK(clk), .Q(sa13[7]) );
  DFFQX1TS \sa23_reg[7]  ( .D(N55), .CK(clk), .Q(sa23[7]) );
  DFFQX1TS \dcnt_reg[0]  ( .D(n988), .CK(clk), .Q(dcnt[0]) );
  DFFXLTS ld_r_reg ( .D(n10366), .CK(clk), .Q(n12765), .QN(n9038) );
  DFFXLTS \dcnt_reg[2]  ( .D(n985), .CK(clk), .QN(n133) );
  AOI211X1TS U1124 ( .A0(n1260), .A1(n139), .B0(n12608), .C0(n12654), .Y(n1262) );
  NOR3BX1TS U1126 ( .AN(n133), .B(dcnt[0]), .C(dcnt[1]), .Y(n1260) );
  OAI2BB2XLTS U1128 ( .B0(text_in_r[35]), .B1(n9470), .A0N(n9469), .A1N(
        text_in_r[35]), .Y(n1268) );
  XOR2X1TS U1129 ( .A(n1269), .B(n1270), .Y(n1266) );
  XOR2X1TS U1130 ( .A(n12662), .B(n1272), .Y(n1270) );
  XNOR2X1TS U1133 ( .A(w2[2]), .B(n1280), .Y(N98) );
  OAI2BB2XLTS U1134 ( .B0(text_in_r[34]), .B1(n12700), .A0N(n1281), .A1N(
        n12716), .Y(n1280) );
  AOI2BB2X1TS U1135 ( .B0(n1282), .B1(n1283), .A0N(n1282), .A1N(n1283), .Y(
        n1281) );
  OAI2BB2XLTS U1138 ( .B0(text_in_r[33]), .B1(n9466), .A0N(n9465), .A1N(
        text_in_r[33]), .Y(n1289) );
  XOR2X1TS U1139 ( .A(n1290), .B(n1291), .Y(n1288) );
  XOR2X1TS U1140 ( .A(n12663), .B(n1293), .Y(n1291) );
  XNOR2X1TS U1143 ( .A(w2[0]), .B(n1299), .Y(N96) );
  OAI2BB2XLTS U1144 ( .B0(text_in_r[32]), .B1(n12710), .A0N(n1300), .A1N(
        n12717), .Y(n1299) );
  AOI2BB2X1TS U1145 ( .B0(n1276), .B1(n1301), .A0N(n1276), .A1N(n1301), .Y(
        n1300) );
  OAI2BB2XLTS U1148 ( .B0(text_in_r[31]), .B1(n9621), .A0N(n9620), .A1N(
        text_in_r[31]), .Y(n1307) );
  XOR2X1TS U1149 ( .A(n1308), .B(n1309), .Y(n1306) );
  XNOR2X1TS U1150 ( .A(n1310), .B(n1311), .Y(n1309) );
  OAI2BB2XLTS U1154 ( .B0(text_in_r[30]), .B1(n9616), .A0N(n9615), .A1N(
        text_in_r[30]), .Y(n1320) );
  XOR2X1TS U1155 ( .A(n1321), .B(n1322), .Y(n1319) );
  XOR2X1TS U1156 ( .A(n1323), .B(n1324), .Y(n1322) );
  OAI2BB2XLTS U1160 ( .B0(text_in_r[29]), .B1(n9611), .A0N(n9610), .A1N(
        text_in_r[29]), .Y(n1333) );
  XOR2X1TS U1161 ( .A(n1334), .B(n1335), .Y(n1332) );
  XOR2X1TS U1162 ( .A(n12660), .B(n1337), .Y(n1335) );
  OAI2BB2XLTS U1166 ( .B0(text_in_r[28]), .B1(n9606), .A0N(n9605), .A1N(
        text_in_r[28]), .Y(n1346) );
  XOR2X1TS U1167 ( .A(n1347), .B(n1348), .Y(n1345) );
  XOR2X1TS U1168 ( .A(n1349), .B(n1350), .Y(n1348) );
  OAI2BB2XLTS U1173 ( .B0(text_in_r[27]), .B1(n9601), .A0N(n9600), .A1N(
        text_in_r[27]), .Y(n1363) );
  XOR2X1TS U1174 ( .A(n1364), .B(n1365), .Y(n1362) );
  XOR2X1TS U1175 ( .A(n1366), .B(n1367), .Y(n1365) );
  AOI2BB2X1TS U1178 ( .B0(n1375), .B1(n9777), .A0N(n9777), .A1N(n1375), .Y(
        n1364) );
  OAI2BB2XLTS U1180 ( .B0(text_in_r[26]), .B1(n9596), .A0N(n9595), .A1N(
        text_in_r[26]), .Y(n1377) );
  XOR2X1TS U1181 ( .A(n1378), .B(n1379), .Y(n1376) );
  XOR2X1TS U1182 ( .A(n1380), .B(n1381), .Y(n1379) );
  OAI2BB2XLTS U1186 ( .B0(text_in_r[25]), .B1(n9592), .A0N(n9591), .A1N(
        text_in_r[25]), .Y(n1390) );
  XOR2X1TS U1187 ( .A(n1391), .B(n1392), .Y(n1389) );
  XOR2X1TS U1188 ( .A(n1393), .B(n1394), .Y(n1392) );
  AOI2BB2X1TS U1191 ( .B0(n12677), .B1(n9234), .A0N(n12677), .A1N(n9234), .Y(
        n1391) );
  XNOR2X1TS U1192 ( .A(w3[24]), .B(n1403), .Y(N80) );
  OAI2BB2XLTS U1193 ( .B0(text_in_r[24]), .B1(n12698), .A0N(n1404), .A1N(
        n12720), .Y(n1403) );
  AOI2BB2X1TS U1194 ( .B0(n1405), .B1(n1406), .A0N(n1405), .A1N(n1406), .Y(
        n1404) );
  XNOR2X1TS U1196 ( .A(w3[23]), .B(n1409), .Y(N71) );
  OAI2BB2XLTS U1197 ( .B0(text_in_r[23]), .B1(n12696), .A0N(n1410), .A1N(
        n12721), .Y(n1409) );
  XNOR2X1TS U1200 ( .A(w3[22]), .B(n1414), .Y(N70) );
  OAI2BB2XLTS U1201 ( .B0(text_in_r[22]), .B1(n12697), .A0N(n1415), .A1N(
        n12722), .Y(n1414) );
  AOI2BB2X1TS U1202 ( .B0(n1336), .B1(n1416), .A0N(n1336), .A1N(n1416), .Y(
        n1415) );
  XNOR2X1TS U1204 ( .A(w3[21]), .B(n1421), .Y(N69) );
  OAI2BB2XLTS U1205 ( .B0(text_in_r[21]), .B1(n12698), .A0N(n1422), .A1N(
        n12724), .Y(n1421) );
  AOI2BB2X1TS U1206 ( .B0(n1359), .B1(n1423), .A0N(n1359), .A1N(n1423), .Y(
        n1422) );
  OAI2BB2XLTS U1209 ( .B0(text_in_r[20]), .B1(n9588), .A0N(n9587), .A1N(
        text_in_r[20]), .Y(n1429) );
  XOR2X1TS U1210 ( .A(n1430), .B(n1431), .Y(n1428) );
  XOR2X1TS U1211 ( .A(n1432), .B(n1375), .Y(n1431) );
  OAI2BB2XLTS U1215 ( .B0(text_in_r[19]), .B1(n9584), .A0N(n9583), .A1N(
        text_in_r[19]), .Y(n1441) );
  XOR2X1TS U1216 ( .A(n1442), .B(n1443), .Y(n1440) );
  XOR2X1TS U1217 ( .A(n1380), .B(n1444), .Y(n1443) );
  XNOR2X1TS U1220 ( .A(w3[18]), .B(n1450), .Y(N66) );
  OAI2BB2XLTS U1221 ( .B0(text_in_r[18]), .B1(n12702), .A0N(n1451), .A1N(
        n12725), .Y(n1450) );
  AOI2BB2X1TS U1222 ( .B0(n9235), .B1(n1452), .A0N(n9234), .A1N(n1452), .Y(
        n1451) );
  OAI2BB2XLTS U1225 ( .B0(text_in_r[17]), .B1(n9579), .A0N(n9578), .A1N(
        text_in_r[17]), .Y(n1458) );
  XOR2X1TS U1226 ( .A(n1459), .B(n1460), .Y(n1457) );
  XOR2X1TS U1227 ( .A(n1405), .B(n1461), .Y(n1460) );
  XNOR2X1TS U1230 ( .A(w3[16]), .B(n1467), .Y(N64) );
  OAI2BB2XLTS U1231 ( .B0(text_in_r[16]), .B1(n12705), .A0N(n1468), .A1N(
        n12727), .Y(n1467) );
  AOI2BB2X1TS U1232 ( .B0(n1438), .B1(n1469), .A0N(n1438), .A1N(n1469), .Y(
        n1468) );
  XNOR2X1TS U1236 ( .A(w3[15]), .B(n1476), .Y(N55) );
  OAI2BB2XLTS U1237 ( .B0(text_in_r[15]), .B1(n12706), .A0N(n1477), .A1N(
        n12728), .Y(n1476) );
  AOI2BB2X1TS U1238 ( .B0(n1478), .B1(n1479), .A0N(n1478), .A1N(n1479), .Y(
        n1477) );
  XNOR2X1TS U1241 ( .A(w3[14]), .B(n1482), .Y(N54) );
  OAI2BB2XLTS U1242 ( .B0(text_in_r[14]), .B1(n12709), .A0N(n1483), .A1N(
        n12729), .Y(n1482) );
  XNOR2X1TS U1246 ( .A(w3[13]), .B(n1487), .Y(N53) );
  OAI2BB2XLTS U1247 ( .B0(text_in_r[13]), .B1(n12706), .A0N(n1488), .A1N(
        n12730), .Y(n1487) );
  AOI2BB2X1TS U1248 ( .B0(n1425), .B1(n1489), .A0N(n1425), .A1N(n1489), .Y(
        n1488) );
  XNOR2X1TS U1249 ( .A(n1435), .B(n1490), .Y(n1489) );
  OAI2BB2XLTS U1253 ( .B0(text_in_r[12]), .B1(n9574), .A0N(n9573), .A1N(
        text_in_r[12]), .Y(n1492) );
  XOR2X1TS U1254 ( .A(n1493), .B(n1494), .Y(n1491) );
  XOR2X1TS U1255 ( .A(n1495), .B(n1496), .Y(n1494) );
  OAI2BB2XLTS U1260 ( .B0(text_in_r[11]), .B1(n9569), .A0N(n9568), .A1N(
        text_in_r[11]), .Y(n1499) );
  XOR2X1TS U1261 ( .A(n1500), .B(n1501), .Y(n1498) );
  XOR2X1TS U1262 ( .A(n1502), .B(n1503), .Y(n1501) );
  AOI2BB2X1TS U1268 ( .B0(w3[0]), .B1(n1408), .A0N(n1408), .A1N(w3[0]), .Y(
        N503) );
  AOI2BB2X1TS U1270 ( .B0(w3[2]), .B1(n9242), .A0N(n9243), .A1N(w3[2]), .Y(
        N501) );
  AOI2BB2X1TS U1271 ( .B0(n9554), .B1(n9246), .A0N(n9247), .A1N(n9554), .Y(
        N500) );
  XNOR2X1TS U1272 ( .A(w3[10]), .B(n1506), .Y(N50) );
  OAI2BB2XLTS U1273 ( .B0(text_in_r[10]), .B1(n12713), .A0N(n1507), .A1N(
        n12732), .Y(n1506) );
  AOI2BB2X1TS U1274 ( .B0(n1454), .B1(n1508), .A0N(n1454), .A1N(n1508), .Y(
        n1507) );
  XNOR2X1TS U1275 ( .A(n1462), .B(n1509), .Y(n1508) );
  AOI2BB2X1TS U1278 ( .B0(w3[5]), .B1(n9254), .A0N(n9255), .A1N(w3[5]), .Y(
        N498) );
  AOI2BB2X1TS U1279 ( .B0(w3[6]), .B1(n9261), .A0N(n9262), .A1N(w3[6]), .Y(
        N497) );
  AOI2BB2X1TS U1280 ( .B0(w3[7]), .B1(n9227), .A0N(n9228), .A1N(w3[7]), .Y(
        N496) );
  AOI2BB2X1TS U1281 ( .B0(w2[0]), .B1(n9224), .A0N(n1511), .A1N(w2[0]), .Y(
        N495) );
  AOI2BB2X1TS U1284 ( .B0(w2[2]), .B1(n9219), .A0N(n9220), .A1N(w2[2]), .Y(
        N493) );
  AOI2BB2X1TS U1288 ( .B0(w2[5]), .B1(n9216), .A0N(n9217), .A1N(w2[5]), .Y(
        N490) );
  OAI2BB2XLTS U1290 ( .B0(text_in_r[9]), .B1(n9564), .A0N(n9563), .A1N(
        text_in_r[9]), .Y(n1522) );
  XOR2X1TS U1291 ( .A(n1523), .B(n1524), .Y(n1521) );
  XOR2X1TS U1292 ( .A(n1525), .B(n1526), .Y(n1524) );
  AOI2BB2X1TS U1297 ( .B0(w2[6]), .B1(n1528), .A0N(n1528), .A1N(w2[6]), .Y(
        N489) );
  AOI2BB2X1TS U1298 ( .B0(w2[7]), .B1(n9212), .A0N(n9213), .A1N(w2[7]), .Y(
        N488) );
  AOI2BB2X1TS U1299 ( .B0(w1[0]), .B1(n9209), .A0N(n9210), .A1N(w1[0]), .Y(
        N487) );
  AOI2BB2X1TS U1301 ( .B0(w1[2]), .B1(n1534), .A0N(n1534), .A1N(w1[2]), .Y(
        N485) );
  AOI2BB2X1TS U1302 ( .B0(n9382), .B1(n1535), .A0N(n1535), .A1N(n9383), .Y(
        N484) );
  AOI2BB2X1TS U1304 ( .B0(w1[5]), .B1(n9206), .A0N(n9207), .A1N(w1[5]), .Y(
        N482) );
  AOI2BB2X1TS U1305 ( .B0(w1[6]), .B1(n9203), .A0N(n1540), .A1N(w1[6]), .Y(
        N481) );
  AOI2BB2X1TS U1306 ( .B0(w1[7]), .B1(n9198), .A0N(n9199), .A1N(w1[7]), .Y(
        N480) );
  XNOR2X1TS U1307 ( .A(w3[8]), .B(n1542), .Y(N48) );
  OAI2BB2XLTS U1308 ( .B0(text_in_r[8]), .B1(n12695), .A0N(n1543), .A1N(n12719), .Y(n1542) );
  XNOR2X1TS U1310 ( .A(n1317), .B(n1471), .Y(n1544) );
  AOI2BB2X1TS U1312 ( .B0(w0[0]), .B1(n9194), .A0N(n9195), .A1N(w0[0]), .Y(
        N479) );
  AOI2BB2X1TS U1314 ( .B0(w0[2]), .B1(n1549), .A0N(n1549), .A1N(w0[2]), .Y(
        N477) );
  AOI2BB2X1TS U1315 ( .B0(n9295), .B1(n9191), .A0N(n9192), .A1N(n9296), .Y(
        N476) );
  AOI2BB2X1TS U1317 ( .B0(w0[5]), .B1(n9187), .A0N(n9188), .A1N(w0[5]), .Y(
        N474) );
  AOI2BB2X1TS U1319 ( .B0(w0[7]), .B1(n9184), .A0N(n9185), .A1N(w0[7]), .Y(
        N472) );
  AOI2BB2X1TS U1320 ( .B0(w3[8]), .B1(n1473), .A0N(n1473), .A1N(w3[8]), .Y(
        N471) );
  AOI2BB2X1TS U1324 ( .B0(w3[10]), .B1(n1456), .A0N(n9773), .A1N(w3[10]), .Y(
        N469) );
  AOI2BB2X1TS U1329 ( .B0(w3[13]), .B1(n1427), .A0N(n1427), .A1N(w3[13]), .Y(
        N466) );
  AOI2BB2X1TS U1331 ( .B0(w3[14]), .B1(n1420), .A0N(n1420), .A1N(w3[14]), .Y(
        N465) );
  AOI2BB2X1TS U1333 ( .B0(w3[15]), .B1(n9230), .A0N(n9231), .A1N(w3[15]), .Y(
        N464) );
  AOI2BB2X1TS U1334 ( .B0(w2[8]), .B1(n9181), .A0N(n9182), .A1N(w2[8]), .Y(
        N463) );
  AOI2BB2X1TS U1336 ( .B0(w2[10]), .B1(n9177), .A0N(n9178), .A1N(w2[10]), .Y(
        N461) );
  AOI2BB2X1TS U1340 ( .B0(w2[14]), .B1(n1567), .A0N(n1567), .A1N(w2[14]), .Y(
        N457) );
  AOI2BB2X1TS U1342 ( .B0(w1[8]), .B1(n1569), .A0N(n1569), .A1N(w1[8]), .Y(
        N455) );
  AOI2BB2X1TS U1348 ( .B0(w1[14]), .B1(n9170), .A0N(n9171), .A1N(w1[14]), .Y(
        N449) );
  AOI2BB2X1TS U1349 ( .B0(w1[15]), .B1(n1582), .A0N(n1582), .A1N(w1[15]), .Y(
        N448) );
  AOI2BB2X1TS U1350 ( .B0(w0[8]), .B1(n1583), .A0N(n1583), .A1N(w0[8]), .Y(
        N447) );
  AOI2BB2X1TS U1355 ( .B0(w0[13]), .B1(n10023), .A0N(n10024), .A1N(w0[13]), 
        .Y(N442) );
  AOI2BB2X1TS U1356 ( .B0(w0[14]), .B1(n9163), .A0N(n9164), .A1N(w0[14]), .Y(
        N441) );
  AOI2BB2X1TS U1357 ( .B0(w0[15]), .B1(n1596), .A0N(n1596), .A1N(w0[15]), .Y(
        N440) );
  AOI2BB2X1TS U1358 ( .B0(w3[16]), .B1(n1398), .A0N(n1398), .A1N(w3[16]), .Y(
        N439) );
  AOI2BB2X1TS U1362 ( .B0(w3[18]), .B1(n1370), .A0N(n9251), .A1N(w3[18]), .Y(
        N437) );
  AOI2BB2X1TS U1367 ( .B0(w3[21]), .B1(n9257), .A0N(n9258), .A1N(w3[21]), .Y(
        N434) );
  AOI2BB2X1TS U1368 ( .B0(w3[22]), .B1(n1310), .A0N(n1310), .A1N(w3[22]), .Y(
        N433) );
  AOI2BB2X1TS U1369 ( .B0(w3[23]), .B1(n9265), .A0N(n9266), .A1N(w3[23]), .Y(
        N432) );
  AOI2BB2X1TS U1370 ( .B0(w2[16]), .B1(n1597), .A0N(n9160), .A1N(w2[16]), .Y(
        N431) );
  AOI2BB2X1TS U1372 ( .B0(w2[18]), .B1(n1601), .A0N(n1601), .A1N(w2[18]), .Y(
        N429) );
  AOI2BB2X1TS U1375 ( .B0(w2[21]), .B1(n1608), .A0N(n1608), .A1N(w2[21]), .Y(
        N426) );
  AOI2BB2X1TS U1376 ( .B0(w2[22]), .B1(n9155), .A0N(n9156), .A1N(w2[22]), .Y(
        N425) );
  AOI2BB2X1TS U1378 ( .B0(w1[16]), .B1(n1611), .A0N(n1611), .A1N(w1[16]), .Y(
        N423) );
  AOI2BB2X1TS U1380 ( .B0(w1[18]), .B1(n9769), .A0N(n9768), .A1N(w1[18]), .Y(
        N421) );
  AOI2BB2X1TS U1383 ( .B0(w1[21]), .B1(n12669), .A0N(n12669), .A1N(w1[21]), 
        .Y(N418) );
  AOI2BB2X1TS U1384 ( .B0(w1[22]), .B1(n9145), .A0N(n9146), .A1N(w1[22]), .Y(
        N417) );
  AOI2BB2X1TS U1385 ( .B0(w1[23]), .B1(n9142), .A0N(n9143), .A1N(w1[23]), .Y(
        N416) );
  AOI2BB2X1TS U1386 ( .B0(w0[16]), .B1(n1625), .A0N(n1625), .A1N(w0[16]), .Y(
        N415) );
  AOI2BB2X1TS U1388 ( .B0(w0[18]), .B1(n12668), .A0N(n12668), .A1N(w0[18]), 
        .Y(N413) );
  AOI2BB2X1TS U1391 ( .B0(w0[21]), .B1(n9133), .A0N(n9134), .A1N(w0[21]), .Y(
        N410) );
  AOI2BB2X1TS U1392 ( .B0(w0[22]), .B1(n10019), .A0N(n10020), .A1N(w0[22]), 
        .Y(N409) );
  AOI2BB2X1TS U1393 ( .B0(w0[23]), .B1(n9130), .A0N(n9131), .A1N(w0[23]), .Y(
        N408) );
  AOI2BB2X1TS U1394 ( .B0(w3[24]), .B1(n1401), .A0N(n1401), .A1N(w3[24]), .Y(
        N407) );
  AOI2BB2X1TS U1409 ( .B0(w2[24]), .B1(n9780), .A0N(n9779), .A1N(w2[24]), .Y(
        N399) );
  AOI2BB2X1TS U1411 ( .B0(w2[26]), .B1(n1287), .A0N(n1287), .A1N(w2[26]), .Y(
        N397) );
  AOI2BB2X1TS U1415 ( .B0(w2[30]), .B1(n1645), .A0N(n1645), .A1N(w2[30]), .Y(
        N393) );
  AOI2BB2X1TS U1417 ( .B0(w1[24]), .B1(n1647), .A0N(n1647), .A1N(w1[24]), .Y(
        N391) );
  XNOR2X1TS U1419 ( .A(w3[7]), .B(n1651), .Y(N39) );
  OAI2BB2XLTS U1420 ( .B0(text_in_r[7]), .B1(n12713), .A0N(n1652), .A1N(n12732), .Y(n1651) );
  AOI2BB2X1TS U1421 ( .B0(n12677), .B1(n1653), .A0N(n1358), .A1N(n1653), .Y(
        n1652) );
  XNOR2X1TS U1422 ( .A(n1475), .B(n1419), .Y(n1653) );
  XNOR2X1TS U1424 ( .A(n9273), .B(n1325), .Y(n1418) );
  NOR4XLTS U1440 ( .A(n1698), .B(n1699), .C(n1700), .D(n1701), .Y(n1697) );
  AOI2BB2X1TS U1446 ( .B0(n10299), .B1(n1724), .A0N(n1725), .A1N(n11143), .Y(
        n1722) );
  NOR4XLTS U1453 ( .A(n1736), .B(n1737), .C(n1738), .D(n1739), .Y(n1735) );
  AOI2BB2X1TS U1459 ( .B0(n10295), .B1(n1762), .A0N(n1763), .A1N(n11121), .Y(
        n1760) );
  AOI2BB2X1TS U1462 ( .B0(w1[26]), .B1(n1770), .A0N(n1770), .A1N(w1[26]), .Y(
        N389) );
  AOI2BB2X1TS U1465 ( .B0(w1[29]), .B1(n1777), .A0N(n9753), .A1N(w1[29]), .Y(
        N386) );
  AOI2BB2X1TS U1466 ( .B0(w1[30]), .B1(n1778), .A0N(n1778), .A1N(w1[30]), .Y(
        N385) );
  XNOR2X1TS U1472 ( .A(w3[6]), .B(n1788), .Y(N38) );
  OAI2BB2XLTS U1473 ( .B0(text_in_r[6]), .B1(n12713), .A0N(n1789), .A1N(n12732), .Y(n1788) );
  AOI2BB2X1TS U1474 ( .B0(n1312), .B1(n1790), .A0N(n9274), .A1N(n1790), .Y(
        n1789) );
  XNOR2X1TS U1475 ( .A(n1323), .B(n1426), .Y(n1790) );
  XNOR2X1TS U1476 ( .A(n1328), .B(n1338), .Y(n1426) );
  NAND4X1TS U1490 ( .A(n1694), .B(n1830), .C(n1831), .D(n1832), .Y(n1829) );
  NAND4X1TS U1496 ( .A(n1850), .B(n1851), .C(n1852), .D(n1853), .Y(n1849) );
  NOR4XLTS U1497 ( .A(n1854), .B(n1855), .C(n1856), .D(n1857), .Y(n1853) );
  NAND2X1TS U1505 ( .A(n11148), .B(n1884), .Y(n1724) );
  NAND4X1TS U1520 ( .A(n1913), .B(n1914), .C(n1915), .D(n1916), .Y(n1912) );
  NOR4XLTS U1521 ( .A(n1917), .B(n1918), .C(n1919), .D(n1920), .Y(n1916) );
  NAND2X1TS U1529 ( .A(n11127), .B(n12346), .Y(n1762) );
  AOI2BB2X1TS U1548 ( .B0(w0[29]), .B1(n1996), .A0N(n1996), .A1N(w0[29]), .Y(
        N378) );
  AOI2BB2X1TS U1549 ( .B0(w0[30]), .B1(n9737), .A0N(n9736), .A1N(w0[30]), .Y(
        N377) );
  AOI2BB2X1TS U1550 ( .B0(w0[31]), .B1(n9100), .A0N(n9101), .A1N(w0[31]), .Y(
        N376) );
  XNOR2X1TS U1551 ( .A(w3[5]), .B(n1999), .Y(N37) );
  OAI2BB2XLTS U1552 ( .B0(text_in_r[5]), .B1(n12711), .A0N(n2000), .A1N(n12732), .Y(n1999) );
  AOI2BB2X1TS U1553 ( .B0(n12660), .B1(n2001), .A0N(n1336), .A1N(n2001), .Y(
        n2000) );
  XNOR2X1TS U1554 ( .A(n1328), .B(n1439), .Y(n2001) );
  XNOR2X1TS U1556 ( .A(n1357), .B(n1341), .Y(n1436) );
  NAND2X1TS U1560 ( .A(n12360), .B(n10616), .Y(n1799) );
  NOR4XLTS U1567 ( .A(n2024), .B(n2025), .C(n2026), .D(n2027), .Y(n1684) );
  XNOR2X1TS U1587 ( .A(n9258), .B(n1424), .Y(n1336) );
  NAND2X1TS U1609 ( .A(n11122), .B(n10251), .Y(n2124) );
  OAI2BB2XLTS U1612 ( .B0(text_in_r[4]), .B1(n9559), .A0N(n9558), .A1N(
        text_in_r[4]), .Y(n2128) );
  XOR2X1TS U1613 ( .A(n2129), .B(n2130), .Y(n2127) );
  XNOR2X1TS U1614 ( .A(n1449), .B(n2131), .Y(n2130) );
  NAND4X1TS U1618 ( .A(n2132), .B(n2133), .C(n2134), .D(n2135), .Y(n1344) );
  NAND3X1TS U1626 ( .A(n2155), .B(n2156), .C(n2157), .Y(n1984) );
  XNOR2X1TS U1634 ( .A(n1352), .B(n1372), .Y(n1449) );
  NAND4X1TS U1647 ( .A(n2203), .B(n2204), .C(n2205), .D(n2206), .Y(n1796) );
  NOR4XLTS U1648 ( .A(n2207), .B(n2208), .C(n2209), .D(n2210), .Y(n2206) );
  NAND2X1TS U1661 ( .A(n12557), .B(n9968), .Y(n1806) );
  XNOR2X1TS U1664 ( .A(n1435), .B(n1343), .Y(n1360) );
  NOR4XLTS U1672 ( .A(n2115), .B(n2248), .C(n2249), .D(n2250), .Y(n1743) );
  OAI221XLTS U1676 ( .A0(n10575), .A1(n10256), .B0(n2260), .B1(n10653), .C0(
        n2261), .Y(n2258) );
  NOR4XLTS U1682 ( .A(n2268), .B(n2269), .C(n2270), .D(n2271), .Y(n2266) );
  NAND4X1TS U1691 ( .A(n2282), .B(n2283), .C(n2284), .D(n2285), .Y(n1911) );
  AOI2BB2X1TS U1699 ( .B0(n10556), .B1(n9756), .A0N(n2297), .A1N(n12085), .Y(
        n2282) );
  NOR4XLTS U1707 ( .A(n2089), .B(n2315), .C(n2316), .D(n2317), .Y(n1705) );
  OAI221XLTS U1711 ( .A0(n10548), .A1(n10280), .B0(n2327), .B1(n10666), .C0(
        n2328), .Y(n2325) );
  NOR4XLTS U1717 ( .A(n2335), .B(n2336), .C(n2337), .D(n2338), .Y(n2333) );
  NAND4X1TS U1726 ( .A(n2349), .B(n2350), .C(n2351), .D(n2352), .Y(n1848) );
  AOI2BB2X1TS U1734 ( .B0(n10528), .B1(n9760), .A0N(n2364), .A1N(n12080), .Y(
        n2349) );
  XNOR2X1TS U1740 ( .A(n1354), .B(n1447), .Y(n1375) );
  NAND4X1TS U1743 ( .A(n2373), .B(n2374), .C(n2375), .D(n2376), .Y(n2372) );
  AOI222XLTS U1745 ( .A0(n11147), .A1(n1706), .B0(n11149), .B1(n11900), .C0(
        n10548), .C1(n10650), .Y(n2378) );
  NOR4XLTS U1747 ( .A(n2381), .B(n2315), .C(n2382), .D(n2383), .Y(n2375) );
  OAI33XLTS U1748 ( .A0(n2341), .A1(n9709), .A2(n10211), .B0(n9939), .B1(
        n10672), .B2(n2386), .Y(n2383) );
  NAND4X1TS U1755 ( .A(n2393), .B(n2394), .C(n2395), .D(n2396), .Y(n2371) );
  NAND4X1TS U1756 ( .A(n2397), .B(n2398), .C(n2399), .D(n2400), .Y(n2075) );
  NOR4XLTS U1757 ( .A(n2401), .B(n2402), .C(n2403), .D(n2404), .Y(n2400) );
  OAI2BB2XLTS U1761 ( .B0(n1725), .B1(n10676), .A0N(n2096), .A1N(n11942), .Y(
        n2403) );
  NOR2BX1TS U1762 ( .AN(n10726), .B(n9061), .Y(n2096) );
  NAND4X1TS U1770 ( .A(n2417), .B(n2418), .C(n2419), .D(n2420), .Y(n2416) );
  AOI222XLTS U1772 ( .A0(n11127), .A1(n1744), .B0(n11126), .B1(n11876), .C0(
        n10575), .C1(n10640), .Y(n2422) );
  NOR4XLTS U1774 ( .A(n2425), .B(n2248), .C(n2426), .D(n2427), .Y(n2419) );
  OAI33XLTS U1775 ( .A0(n2274), .A1(n9705), .A2(n10219), .B0(n9935), .B1(
        n10658), .B2(n2430), .Y(n2427) );
  NAND4X1TS U1782 ( .A(n2437), .B(n2438), .C(n2439), .D(n2440), .Y(n2415) );
  NAND4X1TS U1783 ( .A(n2441), .B(n2442), .C(n2443), .D(n2444), .Y(n2101) );
  NOR4XLTS U1784 ( .A(n2445), .B(n2446), .C(n2447), .D(n2448), .Y(n2444) );
  OAI2BB2XLTS U1788 ( .B0(n1763), .B1(n10662), .A0N(n2122), .A1N(n11931), .Y(
        n2447) );
  NOR2BX1TS U1789 ( .AN(n10700), .B(n9054), .Y(n2122) );
  NAND4X1TS U1796 ( .A(n2458), .B(n2459), .C(n2460), .D(n2461), .Y(n1353) );
  NOR4XLTS U1797 ( .A(n2462), .B(n2048), .C(n2463), .D(n2464), .Y(n2461) );
  NAND2X1TS U1800 ( .A(n11036), .B(n12318), .Y(n2058) );
  OAI2BB2XLTS U1801 ( .B0(n2059), .B1(n12116), .A0N(n2055), .A1N(n10196), .Y(
        n2463) );
  NAND4X1TS U1802 ( .A(n2472), .B(n2473), .C(n2474), .D(n2475), .Y(n2048) );
  NOR4XLTS U1803 ( .A(n2476), .B(n2477), .C(n2478), .D(n2479), .Y(n2475) );
  AOI222XLTS U1811 ( .A0(n10514), .A1(n2493), .B0(n11010), .B1(n2151), .C0(
        n10227), .C1(n2494), .Y(n2489) );
  NOR4XLTS U1812 ( .A(n2495), .B(n2496), .C(n2497), .D(n2498), .Y(n2460) );
  NOR4XLTS U1816 ( .A(n2503), .B(n2504), .C(n2505), .D(n2506), .Y(n2459) );
  XNOR2X1TS U1823 ( .A(n1368), .B(n1382), .Y(n1455) );
  NOR4XLTS U1827 ( .A(n2519), .B(n2187), .C(n2520), .D(n2521), .Y(n2516) );
  NOR4XLTS U1829 ( .A(n2523), .B(n2524), .C(n2525), .D(n2526), .Y(n1792) );
  OAI221XLTS U1836 ( .A0(n12557), .A1(n10690), .B0(n1804), .B1(n11638), .C0(
        n2536), .Y(n2187) );
  NAND2X1TS U1840 ( .A(n10180), .B(n11452), .Y(n1683) );
  NAND3X1TS U1847 ( .A(n2547), .B(n2548), .C(n1687), .Y(n2541) );
  NAND2X1TS U1848 ( .A(n11595), .B(n11917), .Y(n1687) );
  OAI33XLTS U1853 ( .A0(n2557), .A1(n2558), .A2(n10175), .B0(n2557), .B1(
        n10000), .B2(n9697), .Y(n2556) );
  AO22X1TS U1854 ( .A0(n10231), .A1(n2221), .B0(n10616), .B1(n2561), .Y(n2555)
         );
  NAND2X1TS U1857 ( .A(n9932), .B(n9928), .Y(n1802) );
  XNOR2X1TS U1858 ( .A(w3[2]), .B(n2565), .Y(N34) );
  OAI2BB2XLTS U1859 ( .B0(text_in_r[2]), .B1(n12710), .A0N(n2566), .A1N(n12731), .Y(n2565) );
  AOI2BB2X1TS U1860 ( .B0(n1380), .B1(n2567), .A0N(n1380), .A1N(n2567), .Y(
        n2566) );
  XNOR2X1TS U1861 ( .A(n1368), .B(n1466), .Y(n2567) );
  XNOR2X1TS U1863 ( .A(n1388), .B(n1396), .Y(n1465) );
  NAND3X1TS U1865 ( .A(n2568), .B(n2006), .C(n2569), .Y(n1397) );
  NOR4XLTS U1866 ( .A(n2570), .B(n2571), .C(n1795), .D(n2572), .Y(n2569) );
  NAND4X1TS U1872 ( .A(n2580), .B(n2581), .C(n2582), .D(n2583), .Y(n2579) );
  NOR4XLTS U1889 ( .A(n2601), .B(n2602), .C(n2603), .D(n2604), .Y(n1654) );
  NAND4X1TS U1895 ( .A(n2608), .B(n2609), .C(n2610), .D(n2522), .Y(n2593) );
  NAND2X1TS U1896 ( .A(n11507), .B(n11954), .Y(n2522) );
  NAND2X1TS U1902 ( .A(n10680), .B(n9748), .Y(n2227) );
  NAND4X1TS U1907 ( .A(n2473), .B(n2620), .C(n2621), .D(n2622), .Y(n1371) );
  NAND4X1TS U1915 ( .A(n2631), .B(n2632), .C(n2633), .D(n2634), .Y(n2043) );
  OAI222X1TS U1917 ( .A0(n2636), .A1(n11062), .B0(n2637), .B1(n11074), .C0(
        n11833), .C1(n11858), .Y(n2635) );
  OAI221XLTS U1935 ( .A0(n11833), .A1(n10508), .B0(n2663), .B1(n9693), .C0(
        n2664), .Y(n2658) );
  XNOR2X1TS U1940 ( .A(n1369), .B(n9773), .Y(n1380) );
  NOR4XLTS U1942 ( .A(n2671), .B(n2672), .C(n2673), .D(n2674), .Y(n2670) );
  NAND2X1TS U1948 ( .A(n10551), .B(n11577), .Y(n1840) );
  NAND2X1TS U1949 ( .A(n11105), .B(n11943), .Y(n2340) );
  NOR4XLTS U1953 ( .A(n2680), .B(n2681), .C(n2682), .D(n2683), .Y(n2081) );
  NOR4XLTS U1967 ( .A(n1834), .B(n2361), .C(n2412), .D(n2691), .Y(n2669) );
  NAND4X1TS U1969 ( .A(n2693), .B(n2694), .C(n2695), .D(n2696), .Y(n2412) );
  NOR4XLTS U1970 ( .A(n2697), .B(n2698), .C(n2699), .D(n2700), .Y(n2696) );
  NOR4XLTS U1984 ( .A(n2704), .B(n2705), .C(n2706), .D(n2707), .Y(n2703) );
  NAND2X1TS U1990 ( .A(n10579), .B(n11566), .Y(n1903) );
  NAND2X1TS U1991 ( .A(n11088), .B(n11931), .Y(n2273) );
  NOR4XLTS U1995 ( .A(n2713), .B(n2714), .C(n2715), .D(n2716), .Y(n2107) );
  NOR4XLTS U2009 ( .A(n1897), .B(n2294), .C(n2456), .D(n2724), .Y(n2702) );
  NAND4X1TS U2011 ( .A(n2726), .B(n2727), .C(n2728), .D(n2729), .Y(n2456) );
  NOR4XLTS U2012 ( .A(n2730), .B(n2731), .C(n2732), .D(n2733), .Y(n2729) );
  OAI2BB2XLTS U2025 ( .B0(text_in_r[1]), .B1(n9550), .A0N(n9549), .A1N(
        text_in_r[1]), .Y(n2736) );
  XOR2X1TS U2026 ( .A(n2737), .B(n2738), .Y(n2735) );
  XOR2X1TS U2027 ( .A(n9235), .B(n2739), .Y(n2738) );
  NOR4XLTS U2033 ( .A(n2047), .B(n2745), .C(n2746), .D(n2747), .Y(n2744) );
  NAND4X1TS U2039 ( .A(n2754), .B(n2755), .C(n2756), .D(n2757), .Y(n2753) );
  NAND2X1TS U2043 ( .A(n11030), .B(n2151), .Y(n2468) );
  NAND2X1TS U2048 ( .A(n10630), .B(n10620), .Y(n2151) );
  NAND2X1TS U2049 ( .A(n11555), .B(n10598), .Y(n2630) );
  NAND2X1TS U2054 ( .A(n2141), .B(n10948), .Y(n2771) );
  NOR4XLTS U2055 ( .A(n2772), .B(n2773), .C(n2774), .D(n2775), .Y(n2770) );
  NAND2X1TS U2069 ( .A(n12111), .B(n11538), .Y(n2512) );
  NOR4XLTS U2074 ( .A(n2231), .B(n2794), .C(n2795), .D(n2796), .Y(n2793) );
  NOR4XLTS U2077 ( .A(n2798), .B(n2799), .C(n2800), .D(n2801), .Y(n1923) );
  OAI2BB2XLTS U2084 ( .B0(n2431), .B1(n1946), .A0N(n9757), .A1N(n11931), .Y(
        n2795) );
  NAND4X1TS U2087 ( .A(n2806), .B(n2807), .C(n2808), .D(n2809), .Y(n2231) );
  NAND4X1TS U2089 ( .A(n2440), .B(n2811), .C(n2812), .D(n2813), .Y(n2810) );
  NAND2X1TS U2102 ( .A(n12125), .B(n11094), .Y(n2816) );
  NAND4BX1TS U2103 ( .AN(n2823), .B(n2824), .C(n2825), .D(n2826), .Y(n1910) );
  NAND2X1TS U2107 ( .A(n12347), .B(n10997), .Y(n2719) );
  OAI221XLTS U2108 ( .A0(n9979), .A1(n11863), .B0(n12467), .B1(n10569), .C0(
        n2829), .Y(n2823) );
  AOI2BB2X1TS U2122 ( .B0(n10200), .B1(n2120), .A0N(n2844), .A1N(n12085), .Y(
        n2806) );
  NAND2X1TS U2123 ( .A(n11864), .B(n11883), .Y(n2120) );
  NOR4XLTS U2124 ( .A(n2102), .B(n2845), .C(n2846), .D(n2847), .Y(n2792) );
  OAI2BB2XLTS U2125 ( .B0(n2246), .B1(n10215), .A0N(n1755), .A1N(n2814), .Y(
        n2847) );
  NAND4X1TS U2131 ( .A(n2850), .B(n2851), .C(n2852), .D(n2853), .Y(n2849) );
  AOI2BB2X1TS U2136 ( .B0(n11924), .B1(n1927), .A0N(n11573), .A1N(n2856), .Y(
        n2850) );
  NAND2X1TS U2137 ( .A(n11465), .B(n11470), .Y(n1927) );
  NAND2X1TS U2143 ( .A(n10993), .B(n11883), .Y(n1937) );
  NAND4X1TS U2148 ( .A(n1830), .B(n1696), .C(n2868), .D(n2869), .Y(n1464) );
  NOR4XLTS U2149 ( .A(n2298), .B(n2870), .C(n2871), .D(n2872), .Y(n2869) );
  NOR4XLTS U2152 ( .A(n2874), .B(n2875), .C(n2876), .D(n2877), .Y(n1860) );
  OAI2BB2XLTS U2159 ( .B0(n2387), .B1(n1883), .A0N(n9761), .A1N(n11943), .Y(
        n2871) );
  NAND4X1TS U2162 ( .A(n2882), .B(n2883), .C(n2884), .D(n2885), .Y(n2298) );
  NAND4X1TS U2164 ( .A(n2396), .B(n2887), .C(n2888), .D(n2889), .Y(n2886) );
  NAND2X1TS U2177 ( .A(n12139), .B(n11110), .Y(n2892) );
  NAND4BX1TS U2178 ( .AN(n2899), .B(n2900), .C(n2901), .D(n2902), .Y(n1847) );
  NAND2X1TS U2182 ( .A(n12354), .B(n10981), .Y(n2686) );
  OAI221XLTS U2183 ( .A0(n9992), .A1(n11887), .B0(n12483), .B1(n10543), .C0(
        n2905), .Y(n2899) );
  AOI2BB2X1TS U2197 ( .B0(n10203), .B1(n2094), .A0N(n2920), .A1N(n12078), .Y(
        n2882) );
  NAND2X1TS U2198 ( .A(n11888), .B(n11907), .Y(n2094) );
  NOR4XLTS U2199 ( .A(n2076), .B(n2921), .C(n2922), .D(n2923), .Y(n2868) );
  OAI2BB2XLTS U2200 ( .B0(n2313), .B1(n10207), .A0N(n10534), .A1N(n2890), .Y(
        n2923) );
  NAND4X1TS U2206 ( .A(n2926), .B(n2927), .C(n2928), .D(n2929), .Y(n2925) );
  AOI2BB2X1TS U2211 ( .B0(n11937), .B1(n1864), .A0N(n11584), .A1N(n2932), .Y(
        n2926) );
  NAND2X1TS U2212 ( .A(n11478), .B(n11482), .Y(n1864) );
  NAND2X1TS U2218 ( .A(n10978), .B(n11907), .Y(n1874) );
  NAND4X1TS U2227 ( .A(n2945), .B(n2181), .C(n2946), .D(n2947), .Y(n2944) );
  NOR4XLTS U2228 ( .A(n2214), .B(n2226), .C(n2948), .D(n2949), .Y(n2947) );
  NAND2X1TS U2239 ( .A(n10012), .B(n10303), .Y(n2561) );
  OAI2BB2XLTS U2242 ( .B0(n2961), .B1(n1686), .A0N(n10679), .A1N(n2023), .Y(
        n2960) );
  NAND2X1TS U2243 ( .A(n10689), .B(n10606), .Y(n2023) );
  NAND2X1TS U2250 ( .A(n10292), .B(n10602), .Y(n2619) );
  NAND2X1TS U2255 ( .A(n2966), .B(n2967), .Y(n2186) );
  NAND2X1TS U2260 ( .A(n12358), .B(n11917), .Y(n2973) );
  NAND4BX1TS U2262 ( .AN(n2975), .B(n2976), .C(n2977), .D(n2583), .Y(n2178) );
  NAND2X1TS U2263 ( .A(n11424), .B(n11919), .Y(n2583) );
  NOR4XLTS U2268 ( .A(n2979), .B(n2980), .C(n2981), .D(n2982), .Y(n1791) );
  NAND2X1TS U2270 ( .A(n10172), .B(n10232), .Y(n2008) );
  NAND2X1TS U2274 ( .A(n10611), .B(n11596), .Y(n2610) );
  OAI33XLTS U2276 ( .A0(n9044), .A1(n9696), .A2(n10956), .B0(n2986), .B1(n9996), .B2(sa32[7]), .Y(n2980) );
  NAND4X1TS U2279 ( .A(n2988), .B(n2989), .C(n2990), .D(n2991), .Y(n2987) );
  NAND2X1TS U2282 ( .A(n11512), .B(n11158), .Y(n2606) );
  NAND2X1TS U2286 ( .A(n9765), .B(n10287), .Y(n2185) );
  NAND2X1TS U2295 ( .A(n9764), .B(n9927), .Y(n2518) );
  NAND3X1TS U2296 ( .A(n3003), .B(n3004), .C(n3005), .Y(n1813) );
  OAI2BB2XLTS U2299 ( .B0(n2607), .B1(n11046), .A0N(n10232), .A1N(n2978), .Y(
        n3006) );
  NAND2X1TS U2303 ( .A(n11508), .B(n11594), .Y(n3011) );
  NOR4XLTS U2304 ( .A(n3012), .B(n3013), .C(n3014), .D(n3015), .Y(n3010) );
  XNOR2X1TS U2312 ( .A(w3[0]), .B(n3016), .Y(N32) );
  OAI2BB2XLTS U2313 ( .B0(text_in_r[0]), .B1(n12713), .A0N(n3017), .A1N(n12731), .Y(n3016) );
  XNOR2X1TS U2315 ( .A(n1405), .B(n9082), .Y(n3018) );
  NAND4X1TS U2318 ( .A(n1959), .B(n2136), .C(n2743), .D(n3019), .Y(n1413) );
  NOR4XLTS U2319 ( .A(n3020), .B(n3021), .C(n2752), .D(n3022), .Y(n3019) );
  NAND2X1TS U2325 ( .A(n12310), .B(n12106), .Y(n2509) );
  NAND4BX1TS U2326 ( .AN(n3027), .B(n3028), .C(n3029), .D(n3030), .Y(n2752) );
  OAI33XLTS U2330 ( .A0(n9856), .A1(n10626), .A2(n2661), .B0(n2508), .B1(
        sa03[6]), .B2(n10524), .Y(n3032) );
  AOI2BB2X1TS U2332 ( .B0(n9689), .B1(n2055), .A0N(n3035), .A1N(n11834), .Y(
        n3034) );
  NAND2X1TS U2333 ( .A(n10187), .B(n10597), .Y(n2055) );
  NAND2X1TS U2338 ( .A(n10523), .B(n12317), .Y(n1961) );
  AOI2BB2X1TS U2341 ( .B0(n12340), .B1(n11028), .A0N(n11554), .A1N(n1964), .Y(
        n3041) );
  OAI2BB2XLTS U2346 ( .B0(n3043), .B1(n9692), .A0N(n11543), .A1N(n2642), .Y(
        n3036) );
  NAND2X1TS U2350 ( .A(n10950), .B(n11440), .Y(n2511) );
  NAND2X1TS U2353 ( .A(n11542), .B(n11562), .Y(n2648) );
  NAND4X1TS U2354 ( .A(n2481), .B(n2053), .C(n3049), .D(n3050), .Y(n3044) );
  NAND2X1TS U2357 ( .A(n12291), .B(n12452), .Y(n2053) );
  NAND2X1TS U2358 ( .A(n12624), .B(n11538), .Y(n2481) );
  NAND4X1TS U2360 ( .A(n2742), .B(n3054), .C(n3055), .D(n3056), .Y(n3053) );
  NAND2X1TS U2363 ( .A(n12316), .B(n11524), .Y(n2491) );
  NAND2X1TS U2365 ( .A(n11852), .B(n10625), .Y(n2470) );
  NAND4X1TS U2368 ( .A(n3061), .B(n3062), .C(n3063), .D(n3064), .Y(n3060) );
  NAND2X1TS U2374 ( .A(n12291), .B(n11069), .Y(n2634) );
  OAI221XLTS U2378 ( .A0(n11833), .A1(n10188), .B0(n11079), .B1(n12099), .C0(
        n3069), .Y(n3068) );
  NAND4X1TS U2387 ( .A(n3077), .B(n3078), .C(n3079), .D(n2655), .Y(n2137) );
  NAND2X1TS U2388 ( .A(n12623), .B(n10195), .Y(n2655) );
  NOR4XLTS U2397 ( .A(n1659), .B(n3085), .C(n2010), .D(n3086), .Y(n3084) );
  OA22X1TS U2400 ( .A0(n9765), .A1(n11590), .B0(n3089), .B1(n11045), .Y(n3087)
         );
  NAND2X1TS U2402 ( .A(n10008), .B(n9959), .Y(n2213) );
  NAND4X1TS U2403 ( .A(n3090), .B(n3091), .C(n3092), .D(n2212), .Y(n2010) );
  NAND2X1TS U2404 ( .A(n11423), .B(n12181), .Y(n2212) );
  NAND2X1TS U2407 ( .A(n11056), .B(n10179), .Y(n1817) );
  NAND2X1TS U2411 ( .A(n10583), .B(n10616), .Y(n2545) );
  NAND2X1TS U2413 ( .A(n12645), .B(n11955), .Y(n3008) );
  NAND2X1TS U2418 ( .A(n12556), .B(n10015), .Y(n2549) );
  NAND4X1TS U2428 ( .A(n2568), .B(n3101), .C(n3102), .D(n3103), .Y(n1659) );
  NOR4XLTS U2429 ( .A(n2002), .B(n2591), .C(n3104), .D(n3105), .Y(n3103) );
  NAND2X1TS U2436 ( .A(n2220), .B(n10008), .Y(n2222) );
  NAND2X1TS U2439 ( .A(n10179), .B(n11513), .Y(n2991) );
  NAND2X1TS U2442 ( .A(n10171), .B(n11912), .Y(n2951) );
  NAND4X1TS U2448 ( .A(n3113), .B(n3114), .C(n3115), .D(n2548), .Y(n2002) );
  NAND2X1TS U2449 ( .A(n11422), .B(n11052), .Y(n2548) );
  AOI2BB2X1TS U2462 ( .B0(n11595), .B1(n2228), .A0N(n2531), .A1N(n10954), .Y(
        n3120) );
  NAND2X1TS U2463 ( .A(n12160), .B(n10685), .Y(n2228) );
  NAND2X1TS U2466 ( .A(n10292), .B(n10956), .Y(n2201) );
  NAND2X1TS U2468 ( .A(n9967), .B(n10176), .Y(n2221) );
  NAND2X1TS U2474 ( .A(n10004), .B(n10955), .Y(n2978) );
  NAND4X1TS U2476 ( .A(n3122), .B(n3123), .C(n3124), .D(n2532), .Y(n3121) );
  NAND2X1TS U2477 ( .A(n10180), .B(n12186), .Y(n2532) );
  AOI222XLTS U2482 ( .A0(n11454), .A1(n3126), .B0(n11056), .B1(n12325), .C0(
        n11051), .C1(n12194), .Y(n3123) );
  AOI222XLTS U2485 ( .A0(n11823), .A1(n3127), .B0(n11821), .B1(n12646), .C0(
        n11057), .C1(n12360), .Y(n3122) );
  NAND2BX1TS U2496 ( .AN(n9733), .B(n9052), .Y(n1686) );
  OA22X1TS U2507 ( .A0(n9764), .A1(n12161), .B0(n10287), .B1(n1670), .Y(n3135)
         );
  NAND2X1TS U2513 ( .A(n9844), .B(n3130), .Y(n1824) );
  NAND2X1TS U2535 ( .A(n11453), .B(n11158), .Y(n3009) );
  NAND2X1TS U2540 ( .A(n9462), .B(n10354), .Y(n3128) );
  NOR2BX1TS U2548 ( .AN(n2996), .B(n9732), .Y(n2611) );
  NAND2X1TS U2549 ( .A(n11947), .B(n10016), .Y(n3000) );
  NAND2X1TS U2561 ( .A(n9097), .B(n10354), .Y(n2986) );
  NAND2X1TS U2582 ( .A(n9848), .B(n2997), .Y(n3125) );
  XNOR2X1TS U2586 ( .A(n1398), .B(n1470), .Y(n1405) );
  NAND2X1TS U2591 ( .A(n11941), .B(n12296), .Y(n2355) );
  NAND2X1TS U2598 ( .A(n10666), .B(n12352), .Y(n2701) );
  NOR4XLTS U2599 ( .A(n2906), .B(n3150), .C(n3151), .D(n3152), .Y(n2080) );
  NAND2X1TS U2601 ( .A(n10264), .B(n11935), .Y(n2919) );
  AOI2BB2X1TS U2602 ( .B0(n1844), .B1(n2890), .A0N(n12174), .A1N(n1868), .Y(
        n3153) );
  NAND2X1TS U2603 ( .A(n12474), .B(n10650), .Y(n2890) );
  NAND4X1TS U2624 ( .A(n3160), .B(n3161), .C(n3162), .D(n2334), .Y(n2402) );
  NAND2X1TS U2625 ( .A(n11106), .B(n11489), .Y(n2334) );
  NAND4X1TS U2636 ( .A(n2079), .B(n3166), .C(n3167), .D(n3168), .Y(n2672) );
  NOR4XLTS U2637 ( .A(n3169), .B(n2401), .C(n3170), .D(n3171), .Y(n3168) );
  NAND2X1TS U2639 ( .A(n10203), .B(n11111), .Y(n1833) );
  NAND4X1TS U2648 ( .A(n3173), .B(n3174), .C(n3175), .D(n2911), .Y(n2401) );
  NAND2X1TS U2649 ( .A(n9983), .B(n11578), .Y(n2911) );
  NAND2X1TS U2653 ( .A(n10527), .B(n11578), .Y(n2902) );
  NAND2X1TS U2654 ( .A(n12144), .B(n10272), .Y(n2879) );
  NAND2X1TS U2665 ( .A(n3179), .B(n3180), .Y(n2389) );
  NAND2X1TS U2671 ( .A(n10284), .B(n9944), .Y(n2943) );
  NOR4XLTS U2684 ( .A(n2936), .B(n2915), .C(n3187), .D(n3188), .Y(n3167) );
  NAND2X1TS U2696 ( .A(n10675), .B(n11619), .Y(n1872) );
  NAND2X1TS U2709 ( .A(n11618), .B(n10275), .Y(n1870) );
  NAND2X1TS U2711 ( .A(n11582), .B(n11625), .Y(n2409) );
  NOR4XLTS U2714 ( .A(n2874), .B(n3193), .C(n3194), .D(n3195), .Y(n2079) );
  NAND2X1TS U2738 ( .A(n11846), .B(n10204), .Y(n2939) );
  NAND2X1TS U2743 ( .A(sa21[3]), .B(n9124), .Y(n3186) );
  NAND2X1TS U2744 ( .A(n12146), .B(n12374), .Y(n2359) );
  NAND2X1TS U2770 ( .A(sa21[0]), .B(n10060), .Y(n3184) );
  NAND2X1TS U2774 ( .A(n2341), .B(n10726), .Y(n3198) );
  NAND2X1TS U2782 ( .A(n10064), .B(n10331), .Y(n3189) );
  NAND2X1TS U2788 ( .A(n11930), .B(n12302), .Y(n2288) );
  NAND2X1TS U2795 ( .A(n10653), .B(n1947), .Y(n2734) );
  NOR4XLTS U2796 ( .A(n2830), .B(n3210), .C(n3211), .D(n3212), .Y(n2106) );
  NAND2X1TS U2798 ( .A(n10240), .B(n11923), .Y(n2843) );
  AOI2BB2X1TS U2799 ( .B0(n12365), .B1(n2814), .A0N(n12166), .A1N(n1931), .Y(
        n3213) );
  NAND2X1TS U2800 ( .A(n12458), .B(n10641), .Y(n2814) );
  NOR4XLTS U2804 ( .A(n3214), .B(n3215), .C(n3216), .D(n3217), .Y(n3204) );
  NAND4X1TS U2821 ( .A(n3220), .B(n3221), .C(n3222), .D(n2267), .Y(n2446) );
  NAND2X1TS U2822 ( .A(n11088), .B(n11495), .Y(n2267) );
  NAND4X1TS U2833 ( .A(n2105), .B(n3226), .C(n3227), .D(n3228), .Y(n2705) );
  NOR4XLTS U2834 ( .A(n3229), .B(n2445), .C(n3230), .D(n3231), .Y(n3228) );
  NAND2X1TS U2836 ( .A(n10199), .B(n11095), .Y(n1896) );
  NAND4X1TS U2845 ( .A(n3233), .B(n3234), .C(n3235), .D(n2835), .Y(n2445) );
  NAND2X1TS U2846 ( .A(n9971), .B(n11566), .Y(n2835) );
  NAND2X1TS U2850 ( .A(n10557), .B(n11567), .Y(n2826) );
  NAND2X1TS U2851 ( .A(n12130), .B(n10247), .Y(n2803) );
  NAND2X1TS U2862 ( .A(n3239), .B(n3240), .Y(n2433) );
  NAND2X1TS U2868 ( .A(n10260), .B(n9948), .Y(n2867) );
  NOR4XLTS U2881 ( .A(n2860), .B(n2839), .C(n3247), .D(n3248), .Y(n3227) );
  NAND2X1TS U2893 ( .A(n10663), .B(n11602), .Y(n1935) );
  NAND2X1TS U2906 ( .A(n11600), .B(n10252), .Y(n1933) );
  NAND2X1TS U2908 ( .A(n11571), .B(n11607), .Y(n2453) );
  NOR4XLTS U2911 ( .A(n2798), .B(n3253), .C(n3254), .D(n3255), .Y(n2105) );
  NAND2X1TS U2935 ( .A(n11840), .B(n10199), .Y(n2863) );
  NAND2X1TS U2940 ( .A(sa10[3]), .B(n9120), .Y(n3246) );
  NAND2X1TS U2941 ( .A(n12131), .B(n12366), .Y(n2292) );
  NAND2X1TS U2967 ( .A(sa10[0]), .B(n10028), .Y(n3244) );
  NAND2X1TS U2971 ( .A(n2274), .B(n10699), .Y(n3258) );
  NAND2X1TS U2979 ( .A(n10032), .B(n10323), .Y(n3249) );
  NAND4X1TS U2981 ( .A(n3263), .B(n2501), .C(n3264), .D(n3265), .Y(n3262) );
  NOR4XLTS U2982 ( .A(n2487), .B(n3266), .C(n2462), .D(n3267), .Y(n3265) );
  NAND2X1TS U2985 ( .A(n12309), .B(n10184), .Y(n3074) );
  NAND2X1TS U2991 ( .A(n11024), .B(n12452), .Y(n2143) );
  AOI2BB2X1TS U2995 ( .B0(n11442), .B1(n2665), .A0N(n11859), .A1N(n2769), .Y(
        n3271) );
  NOR4XLTS U2998 ( .A(n3272), .B(n3273), .C(n3274), .D(n3275), .Y(n3263) );
  NAND4X1TS U3009 ( .A(n3276), .B(n3277), .C(n3278), .D(n3279), .Y(n2063) );
  AOI2BB2X1TS U3013 ( .B0(n12653), .B1(n3058), .A0N(n2776), .A1N(n11835), .Y(
        n3278) );
  NAND4X1TS U3028 ( .A(n3285), .B(n3286), .C(n3287), .D(n3288), .Y(n2624) );
  NOR4XLTS U3029 ( .A(n2502), .B(n3289), .C(n3290), .D(n3291), .Y(n3288) );
  NAND2X1TS U3031 ( .A(n11041), .B(n9091), .Y(n3069) );
  NAND4X1TS U3034 ( .A(n3294), .B(n3295), .C(n2791), .D(n3296), .Y(n2503) );
  NAND2X1TS U3036 ( .A(n12624), .B(n9091), .Y(n2791) );
  NAND2X1TS U3038 ( .A(n11034), .B(n12116), .Y(n2657) );
  NAND2X1TS U3039 ( .A(n10523), .B(n10592), .Y(n3058) );
  NAND2X1TS U3043 ( .A(n11022), .B(n12613), .Y(n3071) );
  NAND2X1TS U3048 ( .A(n11817), .B(n10515), .Y(n3065) );
  NAND2X1TS U3070 ( .A(n11009), .B(n10589), .Y(n2766) );
  NAND2X1TS U3086 ( .A(n2510), .B(n11554), .Y(n3297) );
  NAND2X1TS U3090 ( .A(sa03[4]), .B(n9067), .Y(n2074) );
  NAND2X1TS U3093 ( .A(n3317), .B(n3318), .Y(n2502) );
  NAND2X1TS U3102 ( .A(n10359), .B(n10364), .Y(n3303) );
  NAND2X1TS U3119 ( .A(n9693), .B(n12116), .Y(n3031) );
  NOR2BX1TS U3121 ( .AN(n3322), .B(n9047), .Y(n2061) );
  AOI2BB2X1TS U3148 ( .B0(n11028), .B1(n2642), .A0N(n10597), .A1N(n2761), .Y(
        n3285) );
  NAND2X1TS U3157 ( .A(n2652), .B(n9530), .Y(n2765) );
  NAND2X1TS U3163 ( .A(n10187), .B(n11548), .Y(n2642) );
  NAND2X1TS U3169 ( .A(n9855), .B(n9522), .Y(n3325) );
  XNOR2X1TS U3175 ( .A(w0[31]), .B(n3326), .Y(N279) );
  OAI2BB2XLTS U3176 ( .B0(text_in_r[127]), .B1(n12709), .A0N(n3327), .A1N(
        n12731), .Y(n3326) );
  AOI2BB2X1TS U3178 ( .B0(n10020), .B1(n9737), .A0N(n9737), .A1N(n10020), .Y(
        n3329) );
  XNOR2X1TS U3180 ( .A(w0[30]), .B(n3333), .Y(N278) );
  OAI2BB2XLTS U3181 ( .B0(text_in_r[126]), .B1(n12711), .A0N(n3334), .A1N(
        n12731), .Y(n3333) );
  XNOR2X1TS U3185 ( .A(w0[29]), .B(n3341), .Y(N277) );
  OAI2BB2XLTS U3186 ( .B0(text_in_r[125]), .B1(n12708), .A0N(n3342), .A1N(
        n12730), .Y(n3341) );
  AOI2BB2X1TS U3187 ( .B0(n3343), .B1(n3344), .A0N(n3343), .A1N(n3344), .Y(
        n3342) );
  AOI2BB2X1TS U3188 ( .B0(n9077), .B1(n1993), .A0N(n12659), .A1N(n9077), .Y(
        n3344) );
  OAI2BB2XLTS U3191 ( .B0(text_in_r[124]), .B1(n9342), .A0N(n9341), .A1N(
        text_in_r[124]), .Y(n3348) );
  XOR2X1TS U3192 ( .A(n3349), .B(n3350), .Y(n3347) );
  XOR2X1TS U3193 ( .A(n3351), .B(n3352), .Y(n3350) );
  OAI2BB2XLTS U3199 ( .B0(text_in_r[123]), .B1(n9338), .A0N(n9337), .A1N(
        text_in_r[123]), .Y(n3358) );
  XOR2X1TS U3200 ( .A(n3359), .B(n3360), .Y(n3357) );
  XOR2X1TS U3201 ( .A(n3361), .B(n3362), .Y(n3360) );
  AOI2BB2X1TS U3205 ( .B0(n12676), .B1(n3366), .A0N(n12676), .A1N(n3366), .Y(
        n3359) );
  XNOR2X1TS U3206 ( .A(w0[26]), .B(n3367), .Y(N274) );
  OAI2BB2XLTS U3207 ( .B0(text_in_r[122]), .B1(n12711), .A0N(n3368), .A1N(
        n12730), .Y(n3367) );
  AOI2BB2X1TS U3208 ( .B0(n3369), .B1(n3370), .A0N(n3369), .A1N(n3370), .Y(
        n3368) );
  AOI2BB2X1TS U3209 ( .B0(n1783), .B1(n3371), .A0N(n3371), .A1N(n1783), .Y(
        n3370) );
  OAI2BB2XLTS U3212 ( .B0(text_in_r[121]), .B1(n9333), .A0N(n9332), .A1N(
        text_in_r[121]), .Y(n3374) );
  XOR2X1TS U3213 ( .A(n3375), .B(n3376), .Y(n3373) );
  XOR2X1TS U3214 ( .A(n3377), .B(n3378), .Y(n3376) );
  AOI2BB2X1TS U3219 ( .B0(n12676), .B1(n9088), .A0N(n3353), .A1N(n9088), .Y(
        n3375) );
  XNOR2X1TS U3220 ( .A(w0[24]), .B(n3382), .Y(N272) );
  OAI2BB2XLTS U3221 ( .B0(text_in_r[120]), .B1(n12711), .A0N(n3383), .A1N(
        n12730), .Y(n3382) );
  AOI2BB2X1TS U3222 ( .B0(n3384), .B1(n3385), .A0N(n3384), .A1N(n3385), .Y(
        n3383) );
  XNOR2X1TS U3224 ( .A(w0[23]), .B(n3387), .Y(N263) );
  OAI2BB2XLTS U3225 ( .B0(text_in_r[119]), .B1(n12710), .A0N(n3388), .A1N(
        n12729), .Y(n3387) );
  XNOR2X1TS U3228 ( .A(w0[22]), .B(n3391), .Y(N262) );
  OAI2BB2XLTS U3229 ( .B0(text_in_r[118]), .B1(n12706), .A0N(n3392), .A1N(
        n12729), .Y(n3391) );
  AOI2BB2X1TS U3230 ( .B0(n9077), .B1(n3393), .A0N(n9078), .A1N(n3393), .Y(
        n3392) );
  XNOR2X1TS U3232 ( .A(w0[21]), .B(n3397), .Y(N261) );
  OAI2BB2XLTS U3233 ( .B0(text_in_r[117]), .B1(n12710), .A0N(n3398), .A1N(
        n12729), .Y(n3397) );
  AOI2BB2X1TS U3234 ( .B0(n3354), .B1(n3399), .A0N(n3354), .A1N(n3399), .Y(
        n3398) );
  AOI2BB2X1TS U3235 ( .B0(n3400), .B1(n10024), .A0N(n10024), .A1N(n3400), .Y(
        n3399) );
  OAI2BB2XLTS U3237 ( .B0(text_in_r[116]), .B1(n9329), .A0N(n9328), .A1N(
        text_in_r[116]), .Y(n3402) );
  XOR2X1TS U3238 ( .A(n3403), .B(n3404), .Y(n3401) );
  XOR2X1TS U3239 ( .A(n3366), .B(n3405), .Y(n3404) );
  OAI2BB2XLTS U3244 ( .B0(text_in_r[115]), .B1(n9325), .A0N(n9324), .A1N(
        text_in_r[115]), .Y(n3411) );
  XOR2X1TS U3245 ( .A(n3412), .B(n3413), .Y(n3410) );
  XNOR2X1TS U3246 ( .A(n3371), .B(n3414), .Y(n3413) );
  XNOR2X1TS U3250 ( .A(w0[18]), .B(n3417), .Y(N258) );
  OAI2BB2XLTS U3251 ( .B0(text_in_r[114]), .B1(n12709), .A0N(n3418), .A1N(
        n12728), .Y(n3417) );
  AOI2BB2X1TS U3252 ( .B0(n9089), .B1(n3419), .A0N(n9088), .A1N(n3419), .Y(
        n3418) );
  OAI2BB2XLTS U3255 ( .B0(text_in_r[113]), .B1(n9321), .A0N(n9320), .A1N(
        text_in_r[113]), .Y(n3424) );
  XOR2X1TS U3256 ( .A(n3425), .B(n3426), .Y(n3423) );
  XOR2X1TS U3257 ( .A(n3384), .B(n3427), .Y(n3426) );
  XNOR2X1TS U3261 ( .A(w0[16]), .B(n3430), .Y(N256) );
  OAI2BB2XLTS U3262 ( .B0(text_in_r[112]), .B1(n12708), .A0N(n3431), .A1N(
        n12728), .Y(n3430) );
  AOI2BB2X1TS U3263 ( .B0(n3407), .B1(n3432), .A0N(n3407), .A1N(n3432), .Y(
        n3431) );
  XNOR2X1TS U3267 ( .A(w0[15]), .B(n3437), .Y(N247) );
  OAI2BB2XLTS U3268 ( .B0(text_in_r[111]), .B1(n12708), .A0N(n3438), .A1N(
        n12728), .Y(n3437) );
  AOI2BB2X1TS U3269 ( .B0(n3439), .B1(n3440), .A0N(n3439), .A1N(n3440), .Y(
        n3438) );
  XNOR2X1TS U3273 ( .A(w0[14]), .B(n3442), .Y(N246) );
  OAI2BB2XLTS U3274 ( .B0(text_in_r[110]), .B1(n12707), .A0N(n3443), .A1N(
        n12727), .Y(n3442) );
  AOI2BB2X1TS U3275 ( .B0(n3444), .B1(n3445), .A0N(n3444), .A1N(n3445), .Y(
        n3443) );
  AOI2BB2X1TS U3276 ( .B0(n10019), .B1(n10023), .A0N(n10023), .A1N(n10019), 
        .Y(n3445) );
  XNOR2X1TS U3278 ( .A(w0[13]), .B(n3446), .Y(N245) );
  OAI2BB2XLTS U3279 ( .B0(text_in_r[109]), .B1(n12706), .A0N(n3447), .A1N(
        n12727), .Y(n3446) );
  AOI2BB2X1TS U3280 ( .B0(n3448), .B1(n3449), .A0N(n3448), .A1N(n3449), .Y(
        n3447) );
  XNOR2X1TS U3282 ( .A(n3400), .B(n1591), .Y(n3448) );
  OAI2BB2XLTS U3284 ( .B0(text_in_r[108]), .B1(n9316), .A0N(n9315), .A1N(
        text_in_r[108]), .Y(n3451) );
  XOR2X1TS U3285 ( .A(n3452), .B(n3453), .Y(n3450) );
  XOR2X1TS U3286 ( .A(n3454), .B(n3455), .Y(n3453) );
  OAI2BB2XLTS U3293 ( .B0(text_in_r[107]), .B1(n9311), .A0N(n9310), .A1N(
        text_in_r[107]), .Y(n3457) );
  XOR2X1TS U3294 ( .A(n3458), .B(n3459), .Y(n3456) );
  XOR2X1TS U3295 ( .A(n3460), .B(n3461), .Y(n3459) );
  XNOR2X1TS U3302 ( .A(w0[10]), .B(n3462), .Y(N242) );
  OAI2BB2XLTS U3303 ( .B0(text_in_r[106]), .B1(n12705), .A0N(n3463), .A1N(
        n12727), .Y(n3462) );
  AOI2BB2X1TS U3304 ( .B0(n1584), .B1(n3464), .A0N(n9168), .A1N(n3464), .Y(
        n3463) );
  XNOR2X1TS U3305 ( .A(n3422), .B(n3465), .Y(n3464) );
  OAI2BB2XLTS U3309 ( .B0(text_in_r[105]), .B1(n9306), .A0N(n9305), .A1N(
        text_in_r[105]), .Y(n3467) );
  XOR2X1TS U3310 ( .A(n3468), .B(n3469), .Y(n3466) );
  XOR2X1TS U3311 ( .A(n3470), .B(n3471), .Y(n3469) );
  XNOR2X1TS U3318 ( .A(w0[8]), .B(n3472), .Y(N240) );
  OAI2BB2XLTS U3319 ( .B0(text_in_r[104]), .B1(n12705), .A0N(n3473), .A1N(
        n12726), .Y(n3472) );
  AOI2BB2X1TS U3320 ( .B0(n9084), .B1(n3474), .A0N(n9085), .A1N(n3474), .Y(
        n3473) );
  XNOR2X1TS U3321 ( .A(n3332), .B(n3434), .Y(n3474) );
  XNOR2X1TS U3324 ( .A(w0[7]), .B(n3475), .Y(N231) );
  OAI2BB2XLTS U3325 ( .B0(text_in_r[103]), .B1(n12704), .A0N(n3476), .A1N(
        n12726), .Y(n3475) );
  AOI2BB2X1TS U3326 ( .B0(n9092), .B1(n3477), .A0N(n9093), .A1N(n3477), .Y(
        n3476) );
  XNOR2X1TS U3327 ( .A(n9080), .B(n3395), .Y(n3477) );
  XOR2X1TS U3329 ( .A(n9736), .B(n3340), .Y(n3396) );
  NAND4BX1TS U3331 ( .AN(n3478), .B(n3479), .C(n3480), .D(n3481), .Y(n1555) );
  NOR4XLTS U3332 ( .A(n3482), .B(n3483), .C(n3484), .D(n3485), .Y(n3481) );
  NAND2X1TS U3341 ( .A(n11416), .B(n12593), .Y(n3515) );
  XNOR2X1TS U3366 ( .A(w0[6]), .B(n3598), .Y(N230) );
  OAI2BB2XLTS U3367 ( .B0(text_in_r[102]), .B1(n12704), .A0N(n3599), .A1N(
        n12726), .Y(n3598) );
  AOI2BB2X1TS U3368 ( .B0(n12670), .B1(n3600), .A0N(n3339), .A1N(n3600), .Y(
        n3599) );
  XOR2X1TS U3369 ( .A(n9736), .B(n3400), .Y(n3600) );
  XNOR2X1TS U3370 ( .A(n1996), .B(n9187), .Y(n3400) );
  NOR4XLTS U3374 ( .A(n3608), .B(n3609), .C(n3610), .D(n3611), .Y(n3607) );
  OAI2BB2XLTS U3377 ( .B0(n12547), .B1(n3618), .A0N(n9903), .A1N(n3620), .Y(
        n3609) );
  NAND4X1TS U3380 ( .A(n3628), .B(n3629), .C(n12037), .D(n11804), .Y(n3601) );
  NOR4XLTS U3388 ( .A(n3654), .B(n3655), .C(n3656), .D(n3657), .Y(n3633) );
  XNOR2X1TS U3393 ( .A(n3394), .B(n10019), .Y(n3339) );
  NAND4X1TS U3408 ( .A(n3715), .B(n3716), .C(n3717), .D(n3718), .Y(n3714) );
  NAND4BX1TS U3415 ( .AN(n3732), .B(n3733), .C(n3734), .D(n3735), .Y(n3731) );
  NAND4X1TS U3433 ( .A(n3781), .B(n3782), .C(n3783), .D(n3784), .Y(n3780) );
  NAND4BX1TS U3440 ( .AN(n3798), .B(n3799), .C(n3800), .D(n3801), .Y(n3797) );
  XNOR2X1TS U3443 ( .A(w0[5]), .B(n3806), .Y(N229) );
  OAI2BB2XLTS U3444 ( .B0(text_in_r[101]), .B1(n12703), .A0N(n3807), .A1N(
        n12726), .Y(n3806) );
  XNOR2X1TS U3446 ( .A(n9078), .B(n3409), .Y(n3808) );
  XNOR2X1TS U3447 ( .A(n1553), .B(n1995), .Y(n3409) );
  NOR4XLTS U3492 ( .A(n3906), .B(n3907), .C(n3908), .D(n3909), .Y(n3905) );
  OAI2BB2XLTS U3493 ( .B0(n3910), .B1(n12539), .A0N(n3911), .A1N(n11248), .Y(
        n3909) );
  OAI2BB2XLTS U3495 ( .B0(n3916), .B1(n12532), .A0N(n9118), .A1N(n3918), .Y(
        n3907) );
  NAND2X1TS U3497 ( .A(n10115), .B(n12018), .Y(n3921) );
  NOR4XLTS U3498 ( .A(n3925), .B(n10877), .C(n10414), .D(n3927), .Y(n3919) );
  OAI2BB2XLTS U3501 ( .B0(text_in_r[100]), .B1(n9301), .A0N(n9300), .A1N(
        text_in_r[100]), .Y(n3932) );
  XOR2X1TS U3502 ( .A(n3933), .B(n3934), .Y(n3931) );
  XNOR2X1TS U3503 ( .A(n3416), .B(n3935), .Y(n3934) );
  XNOR2X1TS U3523 ( .A(n1785), .B(n3365), .Y(n3416) );
  NOR4XLTS U3526 ( .A(n3973), .B(n3974), .C(n3975), .D(n3976), .Y(n3972) );
  NOR4XLTS U3528 ( .A(n3980), .B(n3981), .C(n3982), .D(n3983), .Y(n3978) );
  OAI2BB2XLTS U3533 ( .B0(n3613), .B1(n11805), .A0N(n11793), .A1N(n3992), .Y(
        n3973) );
  NOR4XLTS U3540 ( .A(n4003), .B(n4004), .C(n4005), .D(n4006), .Y(n3604) );
  NOR4XLTS U3542 ( .A(n4009), .B(n4010), .C(n4011), .D(n4012), .Y(n4007) );
  AO22X1TS U3549 ( .A0(n4021), .A1(n11267), .B0(n11793), .B1(n4022), .Y(n4018)
         );
  XNOR2X1TS U3552 ( .A(n1591), .B(n1633), .Y(n3355) );
  NOR4XLTS U3557 ( .A(n4033), .B(n4034), .C(n4035), .D(n4036), .Y(n3526) );
  AOI222XLTS U3559 ( .A0(n12253), .A1(n12002), .B0(n12252), .B1(n10495), .C0(
        n12001), .C1(n12438), .Y(n4038) );
  NAND2X1TS U3563 ( .A(n12587), .B(n11751), .Y(n4041) );
  NOR4XLTS U3565 ( .A(n3711), .B(n4045), .C(n4046), .D(n4047), .Y(n4026) );
  NAND4X1TS U3566 ( .A(n3681), .B(n4048), .C(n4049), .D(n4050), .Y(n4047) );
  OA22X1TS U3569 ( .A0(n9667), .A1(n12009), .B0(n3866), .B1(n10837), .Y(n4048)
         );
  AOI222XLTS U3576 ( .A0(n12438), .A1(n10495), .B0(n11326), .B1(n12059), .C0(
        n12223), .C1(n11404), .Y(n4053) );
  NAND4X1TS U3578 ( .A(n4067), .B(n4068), .C(n4069), .D(n4070), .Y(n3711) );
  NOR4XLTS U3590 ( .A(n4089), .B(n4090), .C(n4091), .D(n4092), .Y(n3565) );
  AOI222XLTS U3592 ( .A0(n12230), .A1(n11987), .B0(n12229), .B1(n10477), .C0(
        n11986), .C1(n12421), .Y(n4094) );
  NAND2X1TS U3596 ( .A(n12578), .B(n11732), .Y(n4097) );
  NOR4XLTS U3598 ( .A(n3777), .B(n4101), .C(n4102), .D(n4103), .Y(n4082) );
  NAND4X1TS U3599 ( .A(n3747), .B(n4104), .C(n4105), .D(n4106), .Y(n4103) );
  OA22X1TS U3602 ( .A0(n9663), .A1(n11996), .B0(n3891), .B1(n10809), .Y(n4104)
         );
  AOI222XLTS U3609 ( .A0(n12422), .A1(n10475), .B0(n11278), .B1(n12052), .C0(
        n12214), .C1(n11392), .Y(n4109) );
  NAND4X1TS U3611 ( .A(n4123), .B(n4124), .C(n4125), .D(n4126), .Y(n3777) );
  OAI2BB2XLTS U3620 ( .B0(text_in_r[99]), .B1(n9295), .A0N(n9295), .A1N(
        text_in_r[99]), .Y(n4138) );
  XOR2X1TS U3621 ( .A(n4139), .B(n4140), .Y(n4137) );
  XOR2X1TS U3622 ( .A(n3366), .B(n9296), .Y(n4140) );
  XNOR2X1TS U3623 ( .A(n1590), .B(n9137), .Y(n3366) );
  NAND4X1TS U3625 ( .A(n4144), .B(n4145), .C(n4146), .D(n4147), .Y(n4143) );
  NAND2X1TS U3628 ( .A(n12516), .B(n11230), .Y(n3538) );
  NOR4XLTS U3631 ( .A(n4154), .B(n4155), .C(n4156), .D(n4157), .Y(n4144) );
  OAI2BB2XLTS U3634 ( .B0(n3868), .B1(n12443), .A0N(n10451), .A1N(n3730), .Y(
        n4155) );
  NAND4BX1TS U3636 ( .AN(n4162), .B(n4163), .C(n4164), .D(n4165), .Y(n4142) );
  NAND2X1TS U3638 ( .A(n10135), .B(n12524), .Y(n4042) );
  NAND4X1TS U3653 ( .A(n4188), .B(n4189), .C(n4190), .D(n4191), .Y(n4187) );
  NAND2X1TS U3656 ( .A(n12498), .B(n11224), .Y(n3577) );
  NOR4XLTS U3659 ( .A(n4198), .B(n4199), .C(n4200), .D(n4201), .Y(n4188) );
  OAI2BB2XLTS U3662 ( .B0(n3893), .B1(n12427), .A0N(n3574), .A1N(n3796), .Y(
        n4199) );
  NAND4BX1TS U3664 ( .AN(n4206), .B(n4207), .C(n4208), .D(n4209), .Y(n4186) );
  NAND2X1TS U3666 ( .A(n10128), .B(n12506), .Y(n4098) );
  XOR2X1TS U3679 ( .A(n1785), .B(n4229), .Y(n4139) );
  NOR4XLTS U3696 ( .A(n4248), .B(n4249), .C(n4250), .D(n4251), .Y(n3622) );
  NAND4BX1TS U3697 ( .AN(n4252), .B(n4253), .C(n4254), .D(n4255), .Y(n4251) );
  NOR4XLTS U3702 ( .A(n4263), .B(n4264), .C(n4265), .D(n4266), .Y(n3970) );
  OAI33XLTS U3714 ( .A0(n9657), .A1(n9172), .A2(n12547), .B0(n9656), .B1(n4282), .B2(n10763), .Y(n4274) );
  NAND3X1TS U3719 ( .A(n4284), .B(n4285), .C(n3904), .Y(n1787) );
  NOR4XLTS U3722 ( .A(n4292), .B(n4293), .C(n4294), .D(n4295), .Y(n4290) );
  NOR4XLTS U3730 ( .A(n4308), .B(n4309), .C(n4310), .D(n4311), .Y(n4285) );
  NAND2X1TS U3737 ( .A(n10777), .B(n12573), .Y(n3911) );
  OAI2BB2XLTS U3738 ( .B0(n9937), .B1(n10456), .A0N(n4325), .A1N(n10796), .Y(
        n4309) );
  NOR4XLTS U3740 ( .A(n4327), .B(n4328), .C(n4329), .D(n4330), .Y(n4284) );
  XNOR2X1TS U3744 ( .A(w0[2]), .B(n4336), .Y(N226) );
  OAI2BB2XLTS U3745 ( .B0(text_in_r[98]), .B1(n12703), .A0N(n4337), .A1N(
        n12725), .Y(n4336) );
  XNOR2X1TS U3747 ( .A(n3371), .B(n3428), .Y(n4338) );
  NOR4XLTS U3753 ( .A(n3608), .B(n4345), .C(n4346), .D(n4347), .Y(n4344) );
  NAND4X1TS U3760 ( .A(n4352), .B(n4353), .C(n4354), .D(n4002), .Y(n3478) );
  NAND2X1TS U3761 ( .A(n10379), .B(n12592), .Y(n4002) );
  NAND4X1TS U3771 ( .A(n4359), .B(n4360), .C(n4361), .D(n4362), .Y(n3810) );
  NOR4XLTS U3773 ( .A(n4364), .B(n4365), .C(n4366), .D(n4367), .Y(n4361) );
  NAND2X1TS U3777 ( .A(n11268), .B(n12073), .Y(n4242) );
  NOR4XLTS U3778 ( .A(n4374), .B(n4375), .C(n4376), .D(n4377), .Y(n3489) );
  NAND2X1TS U3791 ( .A(n4348), .B(n10384), .Y(n3987) );
  NAND2X1TS U3792 ( .A(n10502), .B(n10939), .Y(n4348) );
  XOR2X1TS U3796 ( .A(n3420), .B(n1629), .Y(n3371) );
  NAND4X1TS U3797 ( .A(n4171), .B(n3853), .C(n4150), .D(n4387), .Y(n1629) );
  NOR4XLTS U3798 ( .A(n4388), .B(n4389), .C(n4390), .D(n4391), .Y(n4387) );
  NOR4XLTS U3809 ( .A(n4400), .B(n4401), .C(n4402), .D(n4403), .Y(n4150) );
  NAND2X1TS U3813 ( .A(n10833), .B(n11739), .Y(n3698) );
  NOR4XLTS U3817 ( .A(n4406), .B(n4407), .C(n4408), .D(n4409), .Y(n3853) );
  NOR4XLTS U3823 ( .A(n4415), .B(n4416), .C(n4417), .D(n4418), .Y(n4171) );
  OAI33XLTS U3828 ( .A0(n4424), .A1(n12443), .A2(n4425), .B0(n3871), .B1(
        n10394), .B2(n11169), .Y(n4416) );
  NAND4X1TS U3833 ( .A(n4215), .B(n3878), .C(n4194), .D(n4427), .Y(n1587) );
  NOR4XLTS U3834 ( .A(n4428), .B(n4429), .C(n4430), .D(n4431), .Y(n4427) );
  NOR4XLTS U3845 ( .A(n4440), .B(n4441), .C(n4442), .D(n4443), .Y(n4194) );
  NAND2X1TS U3849 ( .A(n10805), .B(n11719), .Y(n3764) );
  NOR4XLTS U3859 ( .A(n4455), .B(n4456), .C(n4457), .D(n4458), .Y(n4215) );
  OAI33XLTS U3864 ( .A0(n4464), .A1(n12429), .A2(n4465), .B0(n3896), .B1(
        n10382), .B2(n11190), .Y(n4456) );
  NAND2X1TS U3877 ( .A(n11250), .B(n11779), .Y(n3661) );
  NOR4XLTS U3881 ( .A(n4486), .B(n4487), .C(n4488), .D(n4489), .Y(n4484) );
  NAND2X1TS U3883 ( .A(n11780), .B(n10808), .Y(n3966) );
  NAND4X1TS U3887 ( .A(n4493), .B(n4494), .C(n4495), .D(n4496), .Y(n3898) );
  NOR4XLTS U3888 ( .A(n4497), .B(n4498), .C(n4499), .D(n4500), .Y(n4495) );
  OA22X1TS U3892 ( .A0(n11381), .A1(n9938), .B0(n10454), .B1(n4503), .Y(n4493)
         );
  OAI33XLTS U3898 ( .A0(n9682), .A1(n4515), .A2(n11715), .B0(n9683), .B1(n4516), .B2(n12532), .Y(n4507) );
  OAI2BB2XLTS U3902 ( .B0(text_in_r[97]), .B1(n9291), .A0N(n9290), .A1N(
        text_in_r[97]), .Y(n4520) );
  XOR2X1TS U3903 ( .A(n4521), .B(n4522), .Y(n4519) );
  XOR2X1TS U3904 ( .A(n9089), .B(n4523), .Y(n4522) );
  NOR4XLTS U3910 ( .A(n3906), .B(n4529), .C(n4530), .D(n4531), .Y(n4528) );
  NOR4XLTS U3918 ( .A(n4537), .B(n4538), .C(n4539), .D(n4540), .Y(n3631) );
  NAND4X1TS U3927 ( .A(n4548), .B(n4549), .C(n4550), .D(n4551), .Y(n3938) );
  NOR4XLTS U3929 ( .A(n4553), .B(n4554), .C(n4555), .D(n4556), .Y(n4550) );
  NAND4X1TS U3932 ( .A(n4562), .B(n4563), .C(n4564), .D(n4565), .Y(n3654) );
  NAND2X1TS U3941 ( .A(n9679), .B(n3927), .Y(n4322) );
  NAND2X1TS U3945 ( .A(n11761), .B(n9670), .Y(n3927) );
  NOR4XLTS U3960 ( .A(n4589), .B(n4590), .C(n4591), .D(n4592), .Y(n3533) );
  OAI221XLTS U3963 ( .A0(n10486), .A1(n12584), .B0(n12446), .B1(n11362), .C0(
        n4594), .Y(n4591) );
  NAND4X1TS U3968 ( .A(n3674), .B(n4596), .C(n4597), .D(n4598), .Y(n4045) );
  NAND4BX1TS U3974 ( .AN(n4606), .B(n4607), .C(n4608), .D(n4609), .Y(n4605) );
  NAND2X1TS U3981 ( .A(n10915), .B(n12001), .Y(n4147) );
  NAND2X1TS U3986 ( .A(n10140), .B(n4177), .Y(n4414) );
  NOR4XLTS U3990 ( .A(n4622), .B(n3548), .C(n4162), .D(n4623), .Y(n4597) );
  NAND4X1TS U3999 ( .A(n4628), .B(n4629), .C(n4630), .D(n4631), .Y(n4627) );
  OA22X1TS U4000 ( .A0(n12010), .A1(n4632), .B0(n3871), .B1(n9668), .Y(n4630)
         );
  NAND2X1TS U4006 ( .A(n12267), .B(n12515), .Y(n4421) );
  NAND2X1TS U4016 ( .A(n10105), .B(n12405), .Y(n3730) );
  NAND2X1TS U4018 ( .A(n10405), .B(n12002), .Y(n3861) );
  NOR4XLTS U4035 ( .A(n4661), .B(n4662), .C(n4663), .D(n4664), .Y(n3572) );
  OAI221XLTS U4038 ( .A0(n10467), .A1(n12577), .B0(n12428), .B1(n11314), .C0(
        n4666), .Y(n4663) );
  NAND4X1TS U4043 ( .A(n3740), .B(n4668), .C(n4669), .D(n4670), .Y(n4101) );
  NAND4BX1TS U4049 ( .AN(n4678), .B(n4679), .C(n4680), .D(n4681), .Y(n4677) );
  NAND2X1TS U4056 ( .A(n10901), .B(n11986), .Y(n4191) );
  NAND2X1TS U4061 ( .A(n10132), .B(n4221), .Y(n4454) );
  NOR4XLTS U4065 ( .A(n4694), .B(n3587), .C(n4206), .D(n4695), .Y(n4669) );
  NAND2X1TS U4072 ( .A(n10817), .B(n12396), .Y(n3887) );
  NAND4X1TS U4074 ( .A(n4700), .B(n4701), .C(n4702), .D(n4703), .Y(n4699) );
  OA22X1TS U4075 ( .A0(n11996), .A1(n4704), .B0(n3896), .B1(n9672), .Y(n4702)
         );
  NAND4X1TS U4080 ( .A(n4710), .B(n4711), .C(n4712), .D(n4461), .Y(n4709) );
  NAND2X1TS U4081 ( .A(n12244), .B(n12499), .Y(n4461) );
  NAND2X1TS U4083 ( .A(n11309), .B(n11725), .Y(n4711) );
  NAND2X1TS U4091 ( .A(n10113), .B(n12396), .Y(n3796) );
  NAND2X1TS U4093 ( .A(n10409), .B(n11985), .Y(n3886) );
  XNOR2X1TS U4101 ( .A(n1780), .B(n9194), .Y(n3435) );
  NAND4X1TS U4104 ( .A(n4724), .B(n4725), .C(n4726), .D(n4727), .Y(n4723) );
  NAND2X1TS U4105 ( .A(n10926), .B(n9917), .Y(n4727) );
  NOR4XLTS U4106 ( .A(n3982), .B(n4728), .C(n4729), .D(n4730), .Y(n4726) );
  NAND2X1TS U4111 ( .A(n10126), .B(n10934), .Y(n4369) );
  NOR4XLTS U4119 ( .A(n4738), .B(n4739), .C(n4740), .D(n4741), .Y(n4724) );
  OAI2BB2XLTS U4123 ( .B0(n3844), .B1(n10794), .A0N(n11418), .A1N(n4383), .Y(
        n4740) );
  OAI2BB2XLTS U4128 ( .B0(n4744), .B1(n12284), .A0N(n10384), .A1N(n3819), .Y(
        n4738) );
  NAND2X1TS U4129 ( .A(n9660), .B(n10504), .Y(n3819) );
  NAND4X1TS U4130 ( .A(n4745), .B(n4746), .C(n4747), .D(n4748), .Y(n4230) );
  NOR4XLTS U4131 ( .A(n4749), .B(n3980), .C(n4750), .D(n4751), .Y(n4748) );
  NAND2X1TS U4134 ( .A(n4755), .B(n4756), .Y(n3981) );
  NAND2X1TS U4143 ( .A(n10160), .B(n10121), .Y(n4370) );
  OAI33XLTS U4146 ( .A0(n4764), .A1(n9661), .A2(n9698), .B0(n9695), .B1(n10107), .B2(sa33[7]), .Y(n4761) );
  NAND4X1TS U4148 ( .A(n4766), .B(n4767), .C(n4768), .D(n4769), .Y(n4009) );
  NAND2X1TS U4160 ( .A(n11220), .B(n10932), .Y(n4777) );
  OAI2BB2XLTS U4162 ( .B0(n4247), .B1(n12275), .A0N(n11810), .A1N(n4780), .Y(
        n4779) );
  NAND2X1TS U4170 ( .A(n12546), .B(n10793), .Y(n4383) );
  NAND2X1TS U4175 ( .A(n10922), .B(n11387), .Y(n3822) );
  NAND4X1TS U4178 ( .A(n4793), .B(n4794), .C(n4795), .D(n4796), .Y(n4792) );
  NAND2X1TS U4182 ( .A(n10107), .B(n9929), .Y(n4379) );
  XNOR2X1TS U4187 ( .A(w0[0]), .B(n4798), .Y(N224) );
  OAI2BB2XLTS U4188 ( .B0(text_in_r[96]), .B1(n12702), .A0N(n4799), .A1N(
        n12725), .Y(n4798) );
  XNOR2X1TS U4190 ( .A(n3384), .B(n9125), .Y(n4800) );
  NOR4XLTS U4198 ( .A(n4808), .B(n4809), .C(n4810), .D(n4811), .Y(n3961) );
  NAND2X1TS U4200 ( .A(n10814), .B(n10396), .Y(n3922) );
  NAND2X1TS U4203 ( .A(n10138), .B(n10802), .Y(n4331) );
  NAND2X1TS U4206 ( .A(n12620), .B(n12031), .Y(n4291) );
  NAND2X1TS U4207 ( .A(n9176), .B(n11701), .Y(n4485) );
  NAND2X1TS U4216 ( .A(n10390), .B(n10876), .Y(n4496) );
  NAND2X1TS U4221 ( .A(n9922), .B(n10143), .Y(n4300) );
  NOR4XLTS U4222 ( .A(n4826), .B(n4827), .C(n4828), .D(n4829), .Y(n4526) );
  AOI2BB2X1TS U4226 ( .B0(n11214), .B1(n9679), .A0N(n11755), .A1N(n3639), .Y(
        n4830) );
  NAND4X1TS U4238 ( .A(n4842), .B(n4843), .C(n4844), .D(n4845), .Y(n3637) );
  NOR4XLTS U4239 ( .A(n4524), .B(n3937), .C(n4846), .D(n4847), .Y(n4845) );
  NAND2X1TS U4242 ( .A(n10783), .B(n12539), .Y(n4324) );
  NAND2X1TS U4245 ( .A(n12572), .B(n11714), .Y(n4306) );
  NAND4X1TS U4268 ( .A(n4869), .B(n4870), .C(n4871), .D(n4872), .Y(n4553) );
  NAND2X1TS U4272 ( .A(n3917), .B(n11757), .Y(n4837) );
  NOR4XLTS U4283 ( .A(n4882), .B(n4883), .C(n4884), .D(n4885), .Y(n3839) );
  NAND2X1TS U4285 ( .A(n10928), .B(n10130), .Y(n3624) );
  NAND2X1TS U4288 ( .A(n10375), .B(n9934), .Y(n3997) );
  NAND2X1TS U4291 ( .A(n11218), .B(n3498), .Y(n4008) );
  NAND2X1TS U4292 ( .A(n11791), .B(n12044), .Y(n4268) );
  NAND2X1TS U4293 ( .A(n9179), .B(n12072), .Y(n4796) );
  NAND2X1TS U4294 ( .A(n12375), .B(n10380), .Y(n4769) );
  NAND2X1TS U4299 ( .A(n11418), .B(n11273), .Y(n4262) );
  NAND2X1TS U4303 ( .A(n10755), .B(n10123), .Y(n4781) );
  NOR4XLTS U4311 ( .A(n4892), .B(n4893), .C(n4894), .D(n4895), .Y(n4341) );
  OA22X1TS U4313 ( .A0(n9169), .A1(n12064), .B0(n3507), .B1(n11803), .Y(n4897)
         );
  NAND4X1TS U4331 ( .A(n4904), .B(n4905), .C(n4906), .D(n4907), .Y(n3482) );
  NOR4XLTS U4332 ( .A(n4339), .B(n3809), .C(n4908), .D(n4909), .Y(n4907) );
  NAND2X1TS U4334 ( .A(n9934), .B(n3989), .Y(n4016) );
  NAND2X1TS U4335 ( .A(n11707), .B(n9913), .Y(n3989) );
  NAND2X1TS U4338 ( .A(n10794), .B(n12065), .Y(n3992) );
  NAND2X1TS U4339 ( .A(n11708), .B(n12283), .Y(n4780) );
  NAND2X1TS U4343 ( .A(n10787), .B(n10764), .Y(n4022) );
  NAND4X1TS U4349 ( .A(n4912), .B(n4913), .C(n4914), .D(n4915), .Y(n3809) );
  NAND2X1TS U4350 ( .A(n10434), .B(n11274), .Y(n4915) );
  NAND2X1TS U4370 ( .A(n10375), .B(n11799), .Y(n4760) );
  NAND2X1TS U4374 ( .A(n10368), .B(n4925), .Y(n3629) );
  NAND4X1TS U4376 ( .A(n4926), .B(n4927), .C(n4928), .D(n4255), .Y(n4924) );
  NAND2X1TS U4377 ( .A(n10129), .B(n10156), .Y(n4255) );
  NAND2X1TS U4379 ( .A(n10433), .B(n10785), .Y(n4928) );
  NAND2X1TS U4402 ( .A(n9660), .B(n10151), .Y(n4021) );
  NAND4X1TS U4404 ( .A(n4934), .B(n4935), .C(n4936), .D(n4937), .Y(n4364) );
  NAND2X1TS U4411 ( .A(n12277), .B(n10939), .Y(n4260) );
  NAND2X1TS U4417 ( .A(n12387), .B(n11803), .Y(n4900) );
  NAND2BX1TS U4442 ( .AN(n10743), .B(sa33[0]), .Y(n4929) );
  NAND2BX1TS U4467 ( .AN(n9884), .B(n10742), .Y(n4764) );
  NAND2X1TS U4475 ( .A(n12251), .B(n9905), .Y(n4631) );
  NOR4XLTS U4477 ( .A(n4949), .B(n4950), .C(n4951), .D(n4952), .Y(n3852) );
  NAND2X1TS U4479 ( .A(n10916), .B(n10855), .Y(n4602) );
  NAND2X1TS U4480 ( .A(n11737), .B(n12525), .Y(n4609) );
  NOR4XLTS U4485 ( .A(n4953), .B(n4954), .C(n4955), .D(n4956), .Y(n4943) );
  OAI2BB2XLTS U4488 ( .B0(n4633), .B1(n10106), .A0N(n4626), .A1N(n11334), .Y(
        n4955) );
  NAND2X1TS U4504 ( .A(n10485), .B(n9669), .Y(n4626) );
  NAND4X1TS U4505 ( .A(n4960), .B(n4961), .C(n4962), .D(n4963), .Y(n4168) );
  AOI2BB2X1TS U4516 ( .B0(n11745), .B1(n4965), .A0N(n11261), .A1N(n4031), .Y(
        n4961) );
  NAND2X1TS U4518 ( .A(n10485), .B(n10489), .Y(n4965) );
  NAND4X1TS U4520 ( .A(n4167), .B(n3859), .C(n4966), .D(n4967), .Y(n4389) );
  NAND2X1TS U4539 ( .A(n11332), .B(n10760), .Y(n3735) );
  NAND2X1TS U4549 ( .A(n10136), .B(n10450), .Y(n3534) );
  NAND2X1TS U4550 ( .A(n12586), .B(n10761), .Y(n4650) );
  NAND2X1TS U4556 ( .A(n11339), .B(n11244), .Y(n3719) );
  NOR4XLTS U4561 ( .A(n4617), .B(n4078), .C(n3732), .D(n4033), .Y(n4181) );
  NAND2X1TS U4581 ( .A(n10394), .B(n10490), .Y(n4179) );
  NAND2X1TS U4586 ( .A(n12268), .B(n10136), .Y(n4635) );
  NAND2X1TS U4589 ( .A(n11358), .B(n11230), .Y(n4077) );
  NAND2X1TS U4594 ( .A(n10856), .B(n12223), .Y(n4603) );
  NAND2X1TS U4628 ( .A(n9828), .B(n9132), .Y(n4980) );
  NAND2X1TS U4642 ( .A(n9351), .B(n4994), .Y(n3871) );
  NAND2X1TS U4648 ( .A(n9358), .B(n9355), .Y(n3863) );
  NAND2X1TS U4655 ( .A(n10052), .B(n10055), .Y(n4993) );
  NAND2X1TS U4663 ( .A(n9348), .B(sa11[0]), .Y(n4986) );
  NAND2X1TS U4670 ( .A(n12230), .B(n9909), .Y(n4703) );
  NOR4XLTS U4672 ( .A(n5007), .B(n5008), .C(n5009), .D(n5010), .Y(n3877) );
  NAND2X1TS U4674 ( .A(n10900), .B(n4119), .Y(n4674) );
  NAND2X1TS U4675 ( .A(n11721), .B(n12506), .Y(n4681) );
  NAND2X1TS U4699 ( .A(n10468), .B(n9671), .Y(n4698) );
  NAND4X1TS U4700 ( .A(n5018), .B(n5019), .C(n5020), .D(n5021), .Y(n4212) );
  AOI2BB2X1TS U4711 ( .B0(n11725), .B1(n5023), .A0N(n11255), .A1N(n4087), .Y(
        n5019) );
  NAND2X1TS U4713 ( .A(n10468), .B(n10471), .Y(n5023) );
  NAND4X1TS U4715 ( .A(n4211), .B(n3884), .C(n5024), .D(n5025), .Y(n4429) );
  NAND2X1TS U4734 ( .A(n11284), .B(n10772), .Y(n3801) );
  NAND2X1TS U4744 ( .A(n10127), .B(n10442), .Y(n3573) );
  NAND2X1TS U4745 ( .A(n4131), .B(n10773), .Y(n4722) );
  NAND2X1TS U4751 ( .A(n11291), .B(n11237), .Y(n3785) );
  NOR4XLTS U4756 ( .A(n4689), .B(n4134), .C(n3798), .D(n4089), .Y(n4225) );
  NAND2X1TS U4781 ( .A(n12244), .B(n10128), .Y(n4707) );
  NAND2X1TS U4784 ( .A(n11310), .B(n11226), .Y(n4133) );
  NAND2X1TS U4823 ( .A(n9840), .B(n9144), .Y(n5038) );
  NAND2X1TS U4837 ( .A(sa22[4]), .B(n5052), .Y(n3896) );
  NAND2X1TS U4843 ( .A(n9458), .B(n9454), .Y(n3888) );
  NAND2X1TS U4850 ( .A(n10080), .B(n10083), .Y(n5051) );
  NAND2X1TS U4858 ( .A(n9447), .B(n9840), .Y(n5044) );
  NOR4XLTS U4861 ( .A(n5062), .B(n5063), .C(n5064), .D(n5065), .Y(n5061) );
  NOR4XLTS U4870 ( .A(n5066), .B(n5067), .C(n5068), .D(n5069), .Y(n3903) );
  NAND2X1TS U4872 ( .A(n10400), .B(n10802), .Y(n4818) );
  NOR4XLTS U4877 ( .A(n3952), .B(n5071), .C(n5072), .D(n5073), .Y(n4286) );
  OAI2BB2XLTS U4882 ( .B0(n3913), .B1(n12539), .A0N(n4568), .A1N(n10401), .Y(
        n5071) );
  NAND2X1TS U4883 ( .A(n10790), .B(n10407), .Y(n4568) );
  NAND2X1TS U4885 ( .A(n10792), .B(n11775), .Y(n4536) );
  NOR4XLTS U4889 ( .A(n3902), .B(n4292), .C(n5083), .D(n5084), .Y(n5082) );
  NAND2X1TS U4891 ( .A(n10400), .B(n10410), .Y(n4875) );
  OAI2BB2XLTS U4895 ( .B0(n4319), .B1(n12571), .A0N(n9098), .A1N(n9690), .Y(
        n5083) );
  NAND2X1TS U4904 ( .A(n10390), .B(n10396), .Y(n4874) );
  NAND2X1TS U4908 ( .A(n10138), .B(n10395), .Y(n4822) );
  NAND2X1TS U4909 ( .A(n12200), .B(n10806), .Y(n4814) );
  NAND2X1TS U4913 ( .A(n10138), .B(n11213), .Y(n4865) );
  NOR4XLTS U4915 ( .A(n5094), .B(n3951), .C(n5095), .D(n5096), .Y(n5093) );
  NAND2X1TS U4917 ( .A(n10147), .B(n11248), .Y(n4559) );
  NAND2X1TS U4931 ( .A(n10859), .B(n9650), .Y(n4819) );
  AOI2BB2X1TS U4935 ( .B0(n9680), .B1(n4502), .A0N(n9922), .A1N(n4573), .Y(
        n5079) );
  NAND2X1TS U4947 ( .A(n12619), .B(n11780), .Y(n4547) );
  OAI2BB2XLTS U4949 ( .B0(n4474), .B1(n11774), .A0N(n4850), .A1N(n11376), .Y(
        n5105) );
  NAND2X1TS U4950 ( .A(n12491), .B(n12022), .Y(n4850) );
  NAND4X1TS U4962 ( .A(n4313), .B(n5107), .C(n5108), .D(n3960), .Y(n5059) );
  NAND2X1TS U4963 ( .A(n10813), .B(n10411), .Y(n3960) );
  NAND2X1TS U4967 ( .A(n10796), .B(n12201), .Y(n4870) );
  NAND2X1TS U4969 ( .A(n11163), .B(n10308), .Y(n5074) );
  NAND2X1TS U4976 ( .A(n4325), .B(n3668), .Y(n4849) );
  NAND2X1TS U4978 ( .A(n12492), .B(n9676), .Y(n4325) );
  AOI2BB2X1TS U4996 ( .B0(n10137), .B1(n4513), .A0N(n12413), .A1N(n4578), .Y(
        n5114) );
  NAND2X1TS U5002 ( .A(n10406), .B(n11775), .Y(n4513) );
  NAND2X1TS U5006 ( .A(n10314), .B(sa00[1]), .Y(n4516) );
  NAND2X1TS U5025 ( .A(n10116), .B(n11780), .Y(n4560) );
  NAND2X1TS U5027 ( .A(n10319), .B(n5116), .Y(n5110) );
  NAND2X1TS U5049 ( .A(n10307), .B(n11163), .Y(n5111) );
  XNOR2X1TS U5053 ( .A(w1[31]), .B(n5118), .Y(N215) );
  OAI2BB2XLTS U5054 ( .B0(text_in_r[95]), .B1(n12702), .A0N(n5119), .A1N(
        n12725), .Y(n5118) );
  XNOR2X1TS U5058 ( .A(w1[30]), .B(n5127), .Y(N214) );
  OAI2BB2XLTS U5059 ( .B0(text_in_r[94]), .B1(n12701), .A0N(n5128), .A1N(
        n12724), .Y(n5127) );
  AOI2BB2X1TS U5060 ( .B0(n5129), .B1(n5130), .A0N(n5129), .A1N(n5130), .Y(
        n5128) );
  AOI2BB2X1TS U5061 ( .B0(n1622), .B1(n1777), .A0N(n9753), .A1N(n1622), .Y(
        n5130) );
  XNOR2X1TS U5063 ( .A(w1[29]), .B(n5134), .Y(N213) );
  OAI2BB2XLTS U5064 ( .B0(text_in_r[93]), .B1(n12701), .A0N(n5135), .A1N(
        n12724), .Y(n5134) );
  AOI2BB2X1TS U5065 ( .B0(n5136), .B1(n5137), .A0N(n5136), .A1N(n5137), .Y(
        n5135) );
  OAI2BB2XLTS U5069 ( .B0(text_in_r[92]), .B1(n9428), .A0N(n9427), .A1N(
        text_in_r[92]), .Y(n5142) );
  XOR2X1TS U5070 ( .A(n5143), .B(n5144), .Y(n5141) );
  XOR2X1TS U5071 ( .A(n5145), .B(n5146), .Y(n5144) );
  OAI2BB2XLTS U5077 ( .B0(text_in_r[91]), .B1(n9423), .A0N(n9422), .A1N(
        text_in_r[91]), .Y(n5152) );
  XOR2X1TS U5078 ( .A(n5153), .B(n5154), .Y(n5151) );
  XOR2X1TS U5079 ( .A(n5155), .B(n5156), .Y(n5154) );
  AOI2BB2X1TS U5083 ( .B0(n5160), .B1(n12675), .A0N(n12675), .A1N(n5160), .Y(
        n5153) );
  XNOR2X1TS U5084 ( .A(w1[26]), .B(n5161), .Y(N210) );
  OAI2BB2XLTS U5085 ( .B0(text_in_r[90]), .B1(n12700), .A0N(n5162), .A1N(
        n12724), .Y(n5161) );
  AOI2BB2X1TS U5086 ( .B0(n5163), .B1(n5164), .A0N(n5163), .A1N(n5164), .Y(
        n5162) );
  AOI2BB2X1TS U5087 ( .B0(n1650), .B1(n5165), .A0N(n5165), .A1N(n1650), .Y(
        n5164) );
  OAI2BB2XLTS U5092 ( .B0(text_in_r[89]), .B1(n9419), .A0N(n9418), .A1N(
        text_in_r[89]), .Y(n5169) );
  XOR2X1TS U5093 ( .A(n5170), .B(n5171), .Y(n5168) );
  XOR2X1TS U5094 ( .A(n5172), .B(n5173), .Y(n5171) );
  XNOR2X1TS U5100 ( .A(w1[24]), .B(n5178), .Y(N208) );
  OAI2BB2XLTS U5101 ( .B0(text_in_r[88]), .B1(n12701), .A0N(n5179), .A1N(
        n12723), .Y(n5178) );
  AOI2BB2X1TS U5102 ( .B0(n5180), .B1(n5181), .A0N(n5180), .A1N(n5181), .Y(
        n5179) );
  XNOR2X1TS U5104 ( .A(w1[23]), .B(n5183), .Y(N199) );
  OAI2BB2XLTS U5105 ( .B0(text_in_r[87]), .B1(n12700), .A0N(n5184), .A1N(
        n12723), .Y(n5183) );
  XNOR2X1TS U5109 ( .A(w1[22]), .B(n5187), .Y(N198) );
  OAI2BB2XLTS U5110 ( .B0(text_in_r[86]), .B1(n12699), .A0N(n5188), .A1N(
        n12723), .Y(n5187) );
  AOI2BB2X1TS U5111 ( .B0(n9264), .B1(n5189), .A0N(n9264), .A1N(n5189), .Y(
        n5188) );
  XNOR2X1TS U5113 ( .A(w1[21]), .B(n5193), .Y(N197) );
  OAI2BB2XLTS U5114 ( .B0(text_in_r[85]), .B1(n12699), .A0N(n5194), .A1N(
        n12723), .Y(n5193) );
  OAI2BB2XLTS U5118 ( .B0(text_in_r[84]), .B1(n9414), .A0N(n9413), .A1N(
        text_in_r[84]), .Y(n5199) );
  XOR2X1TS U5119 ( .A(n5200), .B(n5201), .Y(n5198) );
  XNOR2X1TS U5120 ( .A(n5160), .B(n5202), .Y(n5201) );
  OAI2BB2XLTS U5125 ( .B0(text_in_r[83]), .B1(n9410), .A0N(n9409), .A1N(
        text_in_r[83]), .Y(n5208) );
  XOR2X1TS U5126 ( .A(n5209), .B(n5210), .Y(n5207) );
  XNOR2X1TS U5127 ( .A(n5165), .B(n5211), .Y(n5210) );
  XNOR2X1TS U5131 ( .A(w1[18]), .B(n5214), .Y(N194) );
  OAI2BB2XLTS U5132 ( .B0(text_in_r[82]), .B1(n12699), .A0N(n5215), .A1N(
        n12722), .Y(n5214) );
  AOI2BB2X1TS U5133 ( .B0(n5176), .B1(n5216), .A0N(n5176), .A1N(n5216), .Y(
        n5215) );
  OAI2BB2XLTS U5137 ( .B0(text_in_r[81]), .B1(n9406), .A0N(n9405), .A1N(
        text_in_r[81]), .Y(n5221) );
  XOR2X1TS U5138 ( .A(n5222), .B(n5223), .Y(n5220) );
  XOR2X1TS U5139 ( .A(n5180), .B(n5224), .Y(n5223) );
  XNOR2X1TS U5143 ( .A(w1[16]), .B(n5227), .Y(N192) );
  OAI2BB2XLTS U5144 ( .B0(text_in_r[80]), .B1(n12697), .A0N(n5228), .A1N(
        n12722), .Y(n5227) );
  AOI2BB2X1TS U5145 ( .B0(n5204), .B1(n5229), .A0N(n5204), .A1N(n5229), .Y(
        n5228) );
  XNOR2X1TS U5149 ( .A(w1[15]), .B(n5234), .Y(N183) );
  OAI2BB2XLTS U5150 ( .B0(text_in_r[79]), .B1(n12699), .A0N(n5235), .A1N(
        n12722), .Y(n5234) );
  AOI2BB2X1TS U5151 ( .B0(n5236), .B1(n5237), .A0N(n5236), .A1N(n5237), .Y(
        n5235) );
  XNOR2X1TS U5154 ( .A(w1[14]), .B(n5239), .Y(N182) );
  OAI2BB2XLTS U5155 ( .B0(text_in_r[78]), .B1(n12697), .A0N(n5240), .A1N(
        n12721), .Y(n5239) );
  AOI2BB2X1TS U5156 ( .B0(n5241), .B1(n5242), .A0N(n5241), .A1N(n5242), .Y(
        n5240) );
  XNOR2X1TS U5159 ( .A(w1[13]), .B(n5243), .Y(N181) );
  OAI2BB2XLTS U5160 ( .B0(text_in_r[77]), .B1(n12698), .A0N(n5244), .A1N(
        n12721), .Y(n5243) );
  AOI2BB2X1TS U5161 ( .B0(n9275), .B1(n5245), .A0N(n9276), .A1N(n5245), .Y(
        n5244) );
  XNOR2X1TS U5162 ( .A(n1577), .B(n5246), .Y(n5245) );
  OAI2BB2XLTS U5165 ( .B0(text_in_r[76]), .B1(n9401), .A0N(n9400), .A1N(
        text_in_r[76]), .Y(n5249) );
  XOR2X1TS U5166 ( .A(n5250), .B(n5251), .Y(n5248) );
  XOR2X1TS U5167 ( .A(n5252), .B(n5253), .Y(n5251) );
  OAI2BB2XLTS U5174 ( .B0(text_in_r[75]), .B1(n9396), .A0N(n9395), .A1N(
        text_in_r[75]), .Y(n5255) );
  XOR2X1TS U5175 ( .A(n5256), .B(n5257), .Y(n5254) );
  XOR2X1TS U5176 ( .A(n5258), .B(n5259), .Y(n5257) );
  XNOR2X1TS U5183 ( .A(w1[10]), .B(n5260), .Y(N178) );
  OAI2BB2XLTS U5184 ( .B0(text_in_r[74]), .B1(n12696), .A0N(n5261), .A1N(
        n12721), .Y(n5260) );
  AOI2BB2X1TS U5185 ( .B0(n1570), .B1(n5262), .A0N(n9174), .A1N(n5262), .Y(
        n5261) );
  XNOR2X1TS U5186 ( .A(n5219), .B(n5263), .Y(n5262) );
  OAI2BB2XLTS U5190 ( .B0(text_in_r[73]), .B1(n9391), .A0N(n9390), .A1N(
        text_in_r[73]), .Y(n5265) );
  XOR2X1TS U5191 ( .A(n5266), .B(n5267), .Y(n5264) );
  XOR2X1TS U5192 ( .A(n5268), .B(n5269), .Y(n5267) );
  XNOR2X1TS U5198 ( .A(w1[8]), .B(n5270), .Y(N176) );
  OAI2BB2XLTS U5199 ( .B0(text_in_r[72]), .B1(n12695), .A0N(n5271), .A1N(
        n12720), .Y(n5270) );
  AOI2BB2X1TS U5200 ( .B0(n9271), .B1(n5272), .A0N(n9272), .A1N(n5272), .Y(
        n5271) );
  XNOR2X1TS U5201 ( .A(n5126), .B(n5231), .Y(n5272) );
  XNOR2X1TS U5204 ( .A(w1[7]), .B(n5273), .Y(N167) );
  OAI2BB2XLTS U5205 ( .B0(text_in_r[71]), .B1(n12695), .A0N(n5274), .A1N(
        n12720), .Y(n5273) );
  AOI2BB2X1TS U5206 ( .B0(n9279), .B1(n5275), .A0N(n9280), .A1N(n5275), .Y(
        n5274) );
  XNOR2X1TS U5207 ( .A(n9267), .B(n5192), .Y(n5275) );
  XNOR2X1TS U5209 ( .A(n1778), .B(n5132), .Y(n5191) );
  NOR4XLTS U5212 ( .A(n5280), .B(n5281), .C(n5282), .D(n5283), .Y(n5279) );
  NAND2X1TS U5221 ( .A(n11206), .B(n12575), .Y(n5313) );
  XNOR2X1TS U5224 ( .A(n9116), .B(n9142), .Y(n5150) );
  XNOR2X1TS U5248 ( .A(w1[6]), .B(n5396), .Y(N166) );
  OAI2BB2XLTS U5249 ( .B0(text_in_r[70]), .B1(n12695), .A0N(n5397), .A1N(
        n12720), .Y(n5396) );
  XNOR2X1TS U5251 ( .A(n5133), .B(n9276), .Y(n5398) );
  NOR4XLTS U5256 ( .A(n5406), .B(n5407), .C(n5408), .D(n5409), .Y(n5405) );
  OAI2BB2XLTS U5259 ( .B0(n12495), .B1(n5416), .A0N(n9953), .A1N(n5418), .Y(
        n5407) );
  NAND4X1TS U5262 ( .A(n9287), .B(n5427), .C(n11976), .D(n11690), .Y(n5399) );
  XNOR2X1TS U5263 ( .A(n5190), .B(n5123), .Y(n5133) );
  NOR4XLTS U5266 ( .A(n5432), .B(n5433), .C(n5434), .D(n5435), .Y(n5431) );
  NAND4X1TS U5267 ( .A(n5436), .B(n5437), .C(n5438), .D(n5439), .Y(n5435) );
  NAND4X1TS U5279 ( .A(n5470), .B(n5471), .C(n5472), .D(n5473), .Y(n5469) );
  NAND4BX1TS U5286 ( .AN(n5487), .B(n5488), .C(n5489), .D(n5490), .Y(n5486) );
  NOR4XLTS U5291 ( .A(n5498), .B(n5499), .C(n5500), .D(n5501), .Y(n5497) );
  NAND4X1TS U5292 ( .A(n5502), .B(n5503), .C(n5504), .D(n5505), .Y(n5501) );
  NAND4X1TS U5304 ( .A(n5536), .B(n5537), .C(n5538), .D(n5539), .Y(n5535) );
  NAND4BX1TS U5311 ( .AN(n5553), .B(n5554), .C(n5555), .D(n5556), .Y(n5552) );
  NAND4X1TS U5315 ( .A(n5565), .B(n5566), .C(n5567), .D(n5568), .Y(n5564) );
  NOR4XLTS U5316 ( .A(n5569), .B(n5570), .C(n5571), .D(n5572), .Y(n5568) );
  NAND2X1TS U5324 ( .A(n11717), .B(n12535), .Y(n5598) );
  XNOR2X1TS U5325 ( .A(w1[5]), .B(n5601), .Y(N165) );
  OAI2BB2XLTS U5326 ( .B0(text_in_r[69]), .B1(n12704), .A0N(n5602), .A1N(
        n12719), .Y(n5601) );
  AOI2BB2X1TS U5327 ( .B0(n9263), .B1(n5603), .A0N(n9263), .A1N(n5603), .Y(
        n5602) );
  XNOR2X1TS U5328 ( .A(n9753), .B(n5203), .Y(n5603) );
  XNOR2X1TS U5329 ( .A(n1538), .B(n1774), .Y(n5203) );
  XNOR2X1TS U5359 ( .A(n1580), .B(n1622), .Y(n5139) );
  NAND4X1TS U5376 ( .A(n5713), .B(n5714), .C(n5715), .D(n5716), .Y(n5712) );
  OAI2BB2XLTS U5385 ( .B0(text_in_r[68]), .B1(n9387), .A0N(n9386), .A1N(
        text_in_r[68]), .Y(n5729) );
  XOR2X1TS U5386 ( .A(n5730), .B(n5731), .Y(n5728) );
  XNOR2X1TS U5387 ( .A(n5213), .B(n5732), .Y(n5731) );
  NOR4XLTS U5392 ( .A(n5736), .B(n5737), .C(n5738), .D(n5739), .Y(n5735) );
  NAND4X1TS U5393 ( .A(n5561), .B(n5740), .C(n5741), .D(n5742), .Y(n5739) );
  OA22X1TS U5396 ( .A0(n9711), .A1(n9981), .B0(n9726), .B1(n5746), .Y(n5740)
         );
  AOI2BB2X1TS U5414 ( .B0(n11679), .B1(n5785), .A0N(n11691), .A1N(n5411), .Y(
        n5775) );
  NOR4XLTS U5416 ( .A(n5787), .B(n5788), .C(n5789), .D(n5790), .Y(n5402) );
  NOR4XLTS U5418 ( .A(n5793), .B(n5794), .C(n5795), .D(n5796), .Y(n5791) );
  AO22X1TS U5425 ( .A0(n5807), .A1(n11341), .B0(n11679), .B1(n5808), .Y(n5804)
         );
  NOR4XLTS U5427 ( .A(n5812), .B(n5813), .C(n5814), .D(n5815), .Y(n5810) );
  XNOR2X1TS U5435 ( .A(n1577), .B(n1619), .Y(n5149) );
  NOR4XLTS U5440 ( .A(n5833), .B(n5834), .C(n5835), .D(n5836), .Y(n5324) );
  AOI222XLTS U5442 ( .A0(n12234), .A1(n12035), .B0(n12233), .B1(n10423), .C0(
        n12034), .C1(n12393), .Y(n5838) );
  NAND2X1TS U5446 ( .A(n12583), .B(n11681), .Y(n5841) );
  NOR4XLTS U5448 ( .A(n5466), .B(n5845), .C(n5846), .D(n5847), .Y(n5826) );
  NAND4X1TS U5449 ( .A(n5436), .B(n5848), .C(n5849), .D(n5850), .Y(n5847) );
  OA22X1TS U5452 ( .A0(n9703), .A1(n12028), .B0(n5696), .B1(n10902), .Y(n5848)
         );
  AOI222XLTS U5459 ( .A0(n12394), .A1(n10423), .B0(n11275), .B1(n5349), .C0(
        n12266), .C1(n11209), .Y(n5853) );
  NAND4X1TS U5461 ( .A(n5867), .B(n5868), .C(n5869), .D(n5870), .Y(n5466) );
  NOR4XLTS U5473 ( .A(n5889), .B(n5890), .C(n5891), .D(n5892), .Y(n5363) );
  AOI222XLTS U5475 ( .A0(n12257), .A1(n12049), .B0(n12256), .B1(n10441), .C0(
        n12048), .C1(n12410), .Y(n5894) );
  NAND2X1TS U5479 ( .A(n12591), .B(n11700), .Y(n5897) );
  NOR4XLTS U5481 ( .A(n5532), .B(n5901), .C(n5902), .D(n5903), .Y(n5882) );
  NAND4X1TS U5482 ( .A(n5502), .B(n5904), .C(n5905), .D(n5906), .Y(n5903) );
  OA22X1TS U5485 ( .A0(n9707), .A1(n12041), .B0(n5721), .B1(n10929), .Y(n5904)
         );
  AOI222XLTS U5492 ( .A0(n12410), .A1(n10441), .B0(n11323), .B1(n5388), .C0(
        n12274), .C1(n11221), .Y(n5909) );
  NAND4X1TS U5494 ( .A(n5923), .B(n5924), .C(n5925), .D(n5926), .Y(n5532) );
  OAI2BB2XLTS U5503 ( .B0(text_in_r[67]), .B1(n9382), .A0N(n9382), .A1N(
        text_in_r[67]), .Y(n5938) );
  XOR2X1TS U5504 ( .A(n5939), .B(n5940), .Y(n5937) );
  XNOR2X1TS U5505 ( .A(n5941), .B(n1773), .Y(n5940) );
  NOR4XLTS U5509 ( .A(n5949), .B(n5950), .C(n5951), .D(n5952), .Y(n5948) );
  NAND2X1TS U5514 ( .A(n10975), .B(n12019), .Y(n5670) );
  NAND4X1TS U5516 ( .A(n5963), .B(n5964), .C(n5965), .D(n5966), .Y(n5943) );
  NAND2X1TS U5519 ( .A(n12054), .B(n12432), .Y(n5969) );
  OAI2BB2XLTS U5521 ( .B0(n5973), .B1(n9722), .A0N(n5974), .A1N(n11348), .Y(
        n5942) );
  NAND3X1TS U5522 ( .A(n5975), .B(n5976), .C(n5977), .Y(n5648) );
  NOR4XLTS U5523 ( .A(n5978), .B(n5979), .C(n5980), .D(n5981), .Y(n5976) );
  OA22X1TS U5530 ( .A0(n10225), .A1(n5759), .B0(n5674), .B1(n5582), .Y(n5993)
         );
  NOR4XLTS U5548 ( .A(n6016), .B(n6017), .C(n6018), .D(n6019), .Y(n5420) );
  NAND4BX1TS U5549 ( .AN(n6020), .B(n6021), .C(n6022), .D(n6023), .Y(n6019) );
  NOR4XLTS U5554 ( .A(n6030), .B(n6031), .C(n6032), .D(n6033), .Y(n5817) );
  OAI33XLTS U5566 ( .A0(n9747), .A1(n6048), .A2(n12494), .B0(n9746), .B1(n6049), .B2(n10979), .Y(n6041) );
  XNOR2X1TS U5570 ( .A(n5160), .B(n9383), .Y(n5939) );
  XOR2X1TS U5571 ( .A(n1576), .B(n9149), .Y(n5160) );
  NAND4X1TS U5573 ( .A(n6054), .B(n6055), .C(n6056), .D(n6057), .Y(n6053) );
  NAND2X1TS U5576 ( .A(n12511), .B(n11407), .Y(n5336) );
  NOR4XLTS U5579 ( .A(n6064), .B(n6065), .C(n6066), .D(n6067), .Y(n6054) );
  OAI2BB2XLTS U5582 ( .B0(n5698), .B1(n12384), .A0N(n10458), .A1N(n5485), .Y(
        n6065) );
  NAND4BX1TS U5584 ( .AN(n6072), .B(n6073), .C(n6074), .D(n6075), .Y(n6052) );
  NAND2X1TS U5586 ( .A(n10161), .B(n12504), .Y(n5842) );
  NAND4X1TS U5601 ( .A(n6098), .B(n6099), .C(n6100), .D(n6101), .Y(n6097) );
  NAND2X1TS U5604 ( .A(n12527), .B(n11413), .Y(n5375) );
  NOR4XLTS U5607 ( .A(n6108), .B(n6109), .C(n6110), .D(n6111), .Y(n6098) );
  OAI2BB2XLTS U5610 ( .B0(n5723), .B1(n12400), .A0N(n10466), .A1N(n5551), .Y(
        n6109) );
  NAND4BX1TS U5612 ( .AN(n6116), .B(n6117), .C(n6118), .D(n6119), .Y(n6096) );
  NAND2X1TS U5614 ( .A(n10170), .B(n12520), .Y(n5898) );
  XNOR2X1TS U5627 ( .A(w1[2]), .B(n6139), .Y(N162) );
  OAI2BB2XLTS U5628 ( .B0(text_in_r[66]), .B1(n12704), .A0N(n6140), .A1N(
        n12718), .Y(n6139) );
  XNOR2X1TS U5630 ( .A(n5165), .B(n5225), .Y(n6141) );
  NOR4XLTS U5636 ( .A(n5406), .B(n6148), .C(n6149), .D(n6150), .Y(n6147) );
  NAND4X1TS U5643 ( .A(n6155), .B(n6156), .C(n6157), .D(n5819), .Y(n5276) );
  NAND2X1TS U5644 ( .A(n10562), .B(n12574), .Y(n5819) );
  NAND4X1TS U5654 ( .A(n6163), .B(n6164), .C(n6165), .D(n6166), .Y(n5605) );
  NOR4XLTS U5656 ( .A(n6168), .B(n6169), .C(n6170), .D(n6171), .Y(n6165) );
  NOR4XLTS U5661 ( .A(n6178), .B(n6179), .C(n6180), .D(n6181), .Y(n5287) );
  NAND2X1TS U5674 ( .A(n10824), .B(n10830), .Y(n6151) );
  XOR2X1TS U5678 ( .A(n5217), .B(n9768), .Y(n5165) );
  NOR4XLTS U5680 ( .A(n6191), .B(n6192), .C(n6193), .D(n6194), .Y(n6190) );
  NOR4XLTS U5691 ( .A(n6203), .B(n6204), .C(n6205), .D(n6206), .Y(n6060) );
  NAND2X1TS U5695 ( .A(n10909), .B(n11694), .Y(n5453) );
  NOR4XLTS U5699 ( .A(n6209), .B(n6210), .C(n6211), .D(n6212), .Y(n5683) );
  NOR4XLTS U5705 ( .A(n6218), .B(n6219), .C(n6220), .D(n6221), .Y(n6081) );
  OAI33XLTS U5710 ( .A0(n6227), .A1(n12384), .A2(n6228), .B0(n5701), .B1(
        n10530), .B2(n11185), .Y(n6219) );
  NAND4X1TS U5715 ( .A(n6125), .B(n5708), .C(n6104), .D(n6230), .Y(n1573) );
  NOR4XLTS U5716 ( .A(n6231), .B(n6232), .C(n6233), .D(n6234), .Y(n6230) );
  NOR4XLTS U5727 ( .A(n6243), .B(n6244), .C(n6245), .D(n6246), .Y(n6104) );
  NAND2X1TS U5731 ( .A(n10936), .B(n11712), .Y(n5519) );
  NOR4XLTS U5741 ( .A(n6258), .B(n6259), .C(n6260), .D(n6261), .Y(n6125) );
  OAI33XLTS U5746 ( .A0(n6267), .A1(n12400), .A2(n6268), .B0(n5726), .B1(
        n10540), .B2(n11202), .Y(n6259) );
  NAND4X1TS U5751 ( .A(n6272), .B(n5650), .C(n6273), .D(n6274), .Y(n6271) );
  NAND4X1TS U5757 ( .A(n6282), .B(n6283), .C(n6284), .D(n6285), .Y(n6281) );
  AOI2BB2X1TS U5779 ( .B0(n11716), .B1(n5988), .A0N(n6315), .A1N(n12014), .Y(
        n6312) );
  OAI33XLTS U5780 ( .A0(n9398), .A1(n11734), .A2(n6317), .B0(n9397), .B1(n6318), .B2(n11752), .Y(n6309) );
  NAND3X1TS U5781 ( .A(n10721), .B(n10194), .C(n6319), .Y(n6307) );
  OAI2BB2XLTS U5784 ( .B0(text_in_r[65]), .B1(n9379), .A0N(n9378), .A1N(
        text_in_r[65]), .Y(n6322) );
  XOR2X1TS U5785 ( .A(n6323), .B(n6324), .Y(n6321) );
  XNOR2X1TS U5786 ( .A(n5177), .B(n6325), .Y(n6324) );
  NAND3X1TS U5791 ( .A(n6328), .B(n5664), .C(n6329), .Y(n6327) );
  NOR4XLTS U5792 ( .A(n6330), .B(n6331), .C(n6332), .D(n6333), .Y(n6329) );
  NAND4X1TS U5800 ( .A(n6342), .B(n6343), .C(n6344), .D(n6345), .Y(n5563) );
  NAND2X1TS U5803 ( .A(n11740), .B(n12534), .Y(n5966) );
  NAND4X1TS U5809 ( .A(n6353), .B(n6354), .C(n6355), .D(n6356), .Y(n5737) );
  NOR4XLTS U5811 ( .A(n6357), .B(n6358), .C(n6359), .D(n6360), .Y(n6355) );
  NAND4X1TS U5814 ( .A(n6366), .B(n6367), .C(n6368), .D(n6369), .Y(n5571) );
  NAND2X1TS U5821 ( .A(n12431), .B(n10963), .Y(n6294) );
  NAND2X1TS U5826 ( .A(n10177), .B(n5995), .Y(n5961) );
  NAND2X1TS U5827 ( .A(n10173), .B(n9388), .Y(n5995) );
  XNOR2X1TS U5831 ( .A(n9173), .B(n1614), .Y(n5177) );
  NOR4XLTS U5843 ( .A(n6389), .B(n6390), .C(n6391), .D(n6392), .Y(n5331) );
  OAI221XLTS U5846 ( .A0(n10432), .A1(n9335), .B0(n12385), .B1(n11239), .C0(
        n6394), .Y(n6391) );
  NAND4X1TS U5851 ( .A(n5429), .B(n6396), .C(n6397), .D(n6398), .Y(n5845) );
  NAND4BX1TS U5857 ( .AN(n6406), .B(n6407), .C(n6408), .D(n6409), .Y(n6405) );
  NAND2X1TS U5864 ( .A(n10853), .B(n12034), .Y(n6057) );
  NAND2X1TS U5869 ( .A(n10158), .B(n6087), .Y(n6217) );
  NOR4XLTS U5873 ( .A(n6422), .B(n5346), .C(n6072), .D(n6423), .Y(n6397) );
  NAND2X1TS U5880 ( .A(n10897), .B(n12415), .Y(n5692) );
  NAND4X1TS U5882 ( .A(n6428), .B(n6429), .C(n6430), .D(n6431), .Y(n6427) );
  OA22X1TS U5883 ( .A0(n12028), .A1(n6432), .B0(n5701), .B1(n9770), .Y(n6430)
         );
  NAND4X1TS U5888 ( .A(n6438), .B(n6439), .C(n6440), .D(n6224), .Y(n6437) );
  NAND2X1TS U5889 ( .A(n12217), .B(n12512), .Y(n6224) );
  NAND2X1TS U5891 ( .A(n11246), .B(n11686), .Y(n6439) );
  NAND2X1TS U5899 ( .A(n10209), .B(n12417), .Y(n5485) );
  NAND2X1TS U5901 ( .A(n10582), .B(n12036), .Y(n5691) );
  NOR4XLTS U5918 ( .A(n6461), .B(n6462), .C(n6463), .D(n6464), .Y(n5370) );
  OAI221XLTS U5921 ( .A0(n10449), .A1(n12588), .B0(n12402), .B1(n11287), .C0(
        n6466), .Y(n6463) );
  NAND4X1TS U5926 ( .A(n5495), .B(n6468), .C(n6469), .D(n6470), .Y(n5901) );
  NAND4BX1TS U5932 ( .AN(n6478), .B(n6479), .C(n6480), .D(n6481), .Y(n6477) );
  NAND2X1TS U5939 ( .A(n10868), .B(n12049), .Y(n6101) );
  NAND2X1TS U5944 ( .A(n10166), .B(n6131), .Y(n6257) );
  NOR4XLTS U5948 ( .A(n6494), .B(n5385), .C(n6116), .D(n6495), .Y(n6469) );
  NAND2X1TS U5955 ( .A(n10924), .B(n12423), .Y(n5717) );
  NAND4X1TS U5957 ( .A(n6500), .B(n6501), .C(n6502), .D(n6503), .Y(n6499) );
  OA22X1TS U5958 ( .A0(n12042), .A1(n6504), .B0(n5726), .B1(n9775), .Y(n6502)
         );
  NAND2X1TS U5964 ( .A(n12240), .B(n12528), .Y(n6264) );
  NAND2X1TS U5974 ( .A(n10217), .B(n12425), .Y(n5551) );
  NAND2X1TS U5976 ( .A(n10586), .B(n12050), .Y(n5716) );
  XNOR2X1TS U5984 ( .A(n1647), .B(n9209), .Y(n5232) );
  NAND2X1TS U5994 ( .A(n10242), .B(n10836), .Y(n6173) );
  NAND2X1TS U6009 ( .A(n10413), .B(n11672), .Y(n5779) );
  NAND2X1TS U6012 ( .A(n9758), .B(n10826), .Y(n5614) );
  NAND4X1TS U6013 ( .A(n6545), .B(n6546), .C(n6547), .D(n6548), .Y(n5997) );
  NOR4XLTS U6014 ( .A(n6549), .B(n5812), .C(n6550), .D(n6551), .Y(n6548) );
  NAND2X1TS U6017 ( .A(n6555), .B(n6556), .Y(n5813) );
  NAND2X1TS U6026 ( .A(n10142), .B(n9993), .Y(n6174) );
  OAI33XLTS U6029 ( .A0(n6564), .A1(n9759), .A2(n9789), .B0(n9786), .B1(n10206), .B2(sa30[7]), .Y(n6561) );
  NAND4X1TS U6031 ( .A(n6566), .B(n6567), .C(n6568), .D(n6569), .Y(n5793) );
  NAND2X1TS U6043 ( .A(n11396), .B(n10834), .Y(n6577) );
  OAI2BB2XLTS U6045 ( .B0(n6014), .B1(n12212), .A0N(n11979), .A1N(n6580), .Y(
        n6579) );
  NAND2X1TS U6053 ( .A(n12496), .B(n10957), .Y(n6187) );
  NAND2X1TS U6058 ( .A(n10847), .B(n11672), .Y(n5617) );
  NAND4X1TS U6061 ( .A(n6593), .B(n6594), .C(n6595), .D(n6596), .Y(n6592) );
  NAND2X1TS U6065 ( .A(n10205), .B(n9767), .Y(n6183) );
  XNOR2X1TS U6070 ( .A(w1[0]), .B(n6598), .Y(N160) );
  OAI2BB2XLTS U6071 ( .B0(text_in_r[64]), .B1(n12696), .A0N(n6599), .A1N(
        n12717), .Y(n6598) );
  XNOR2X1TS U6073 ( .A(n5180), .B(n9317), .Y(n6600) );
  NAND4X1TS U6077 ( .A(n6353), .B(n5765), .C(n6604), .D(n6605), .Y(n6603) );
  NAND4X1TS U6081 ( .A(n6610), .B(n6611), .C(n6301), .D(n5985), .Y(n6609) );
  NAND2X1TS U6082 ( .A(n12542), .B(n12535), .Y(n5985) );
  NAND2X1TS U6083 ( .A(n9977), .B(n11998), .Y(n6301) );
  NAND2X1TS U6084 ( .A(n12433), .B(n10942), .Y(n6611) );
  NAND2X1TS U6087 ( .A(n11723), .B(n10577), .Y(n5652) );
  NAND2X1TS U6090 ( .A(n10546), .B(n11331), .Y(n5970) );
  NAND2X1TS U6097 ( .A(n11718), .B(n12063), .Y(n6285) );
  NAND4X1TS U6100 ( .A(n6624), .B(n6625), .C(n6626), .D(n6627), .Y(n6330) );
  NAND2X1TS U6103 ( .A(n11741), .B(n10249), .Y(n6278) );
  AOI2BB2X1TS U6107 ( .B0(n12278), .B1(n10178), .A0N(n12005), .A1N(n5589), .Y(
        n6624) );
  NAND4X1TS U6119 ( .A(n6641), .B(n6642), .C(n6643), .D(n6644), .Y(n5562) );
  NOR4XLTS U6120 ( .A(n6326), .B(n5736), .C(n6645), .D(n6646), .Y(n6644) );
  NAND2X1TS U6123 ( .A(n10474), .B(n12287), .Y(n5962) );
  NAND2X1TS U6126 ( .A(n12020), .B(n11753), .Y(n5988) );
  NAND4X1TS U6148 ( .A(n6667), .B(n6668), .C(n6669), .D(n6670), .Y(n6357) );
  NAND2X1TS U6150 ( .A(n6672), .B(n6673), .Y(n6671) );
  NAND2X1TS U6151 ( .A(n11747), .B(n12006), .Y(n6633) );
  NAND2X1TS U6153 ( .A(n9388), .B(n11992), .Y(n6289) );
  NOR4XLTS U6165 ( .A(n6681), .B(n6682), .C(n6683), .D(n6684), .Y(n5634) );
  NAND2X1TS U6167 ( .A(n10842), .B(n9998), .Y(n5422) );
  NAND2X1TS U6170 ( .A(n10559), .B(n9990), .Y(n5822) );
  NAND4X1TS U6172 ( .A(n6569), .B(n6596), .C(n6035), .D(n5792), .Y(n6682) );
  NAND2X1TS U6173 ( .A(n11395), .B(n9637), .Y(n5792) );
  NAND2X1TS U6174 ( .A(n11677), .B(n11669), .Y(n6035) );
  NAND2X1TS U6175 ( .A(n9375), .B(n11696), .Y(n6596) );
  NAND2X1TS U6176 ( .A(n12447), .B(n10563), .Y(n6569) );
  NAND2X1TS U6181 ( .A(n11206), .B(n11336), .Y(n6029) );
  NAND2X1TS U6185 ( .A(n10990), .B(n10185), .Y(n6581) );
  NOR4XLTS U6193 ( .A(n6691), .B(n6692), .C(n6693), .D(n6694), .Y(n6144) );
  OA22X1TS U6195 ( .A0(n9356), .A1(n12196), .B0(n5305), .B1(n11689), .Y(n6696)
         );
  NAND4X1TS U6213 ( .A(n6703), .B(n6704), .C(n6705), .D(n6706), .Y(n5280) );
  NOR4XLTS U6214 ( .A(n6142), .B(n5604), .C(n6707), .D(n6708), .Y(n6706) );
  NAND2X1TS U6216 ( .A(n9990), .B(n5783), .Y(n5802) );
  NAND2X1TS U6217 ( .A(n11401), .B(n9965), .Y(n5783) );
  NAND2X1TS U6220 ( .A(n10958), .B(n12197), .Y(n5785) );
  NAND2X1TS U6221 ( .A(n11402), .B(n12204), .Y(n6580) );
  NAND2X1TS U6225 ( .A(n10500), .B(n10980), .Y(n5808) );
  NAND4X1TS U6231 ( .A(n6711), .B(n6712), .C(n6713), .D(n6714), .Y(n5604) );
  NAND2X1TS U6232 ( .A(n10492), .B(n11335), .Y(n6714) );
  NAND2X1TS U6252 ( .A(n10559), .B(n11684), .Y(n6560) );
  NAND2X1TS U6256 ( .A(sa30[4]), .B(n6724), .Y(n5427) );
  NAND4X1TS U6258 ( .A(n6725), .B(n6726), .C(n6727), .D(n6023), .Y(n6723) );
  NAND2X1TS U6259 ( .A(n9997), .B(n10146), .Y(n6023) );
  NAND2X1TS U6261 ( .A(n10491), .B(n11378), .Y(n6727) );
  NAND2X1TS U6283 ( .A(n9758), .B(n10149), .Y(n5807) );
  NAND4X1TS U6285 ( .A(n6733), .B(n6734), .C(n6735), .D(n6736), .Y(n6168) );
  NAND2X1TS U6292 ( .A(n12212), .B(n10829), .Y(n6027) );
  NAND2X1TS U6298 ( .A(n12439), .B(n11689), .Y(n6699) );
  NAND2BX1TS U6323 ( .AN(n10710), .B(sa30[0]), .Y(n6728) );
  NAND2BX1TS U6350 ( .AN(n9808), .B(n10710), .Y(n6564) );
  NAND2X1TS U6358 ( .A(n12232), .B(n9957), .Y(n6431) );
  NOR4XLTS U6360 ( .A(n6748), .B(n6749), .C(n6750), .D(n6751), .Y(n5682) );
  NAND2X1TS U6362 ( .A(n10852), .B(n10886), .Y(n6402) );
  NAND2X1TS U6363 ( .A(n11692), .B(n12502), .Y(n6409) );
  NOR4XLTS U6368 ( .A(n6752), .B(n6753), .C(n6754), .D(n6755), .Y(n6742) );
  OAI2BB2XLTS U6371 ( .B0(n6433), .B1(n10210), .A0N(n6426), .A1N(n11271), .Y(
        n6754) );
  NAND2X1TS U6387 ( .A(n10431), .B(n9771), .Y(n6426) );
  NAND4X1TS U6388 ( .A(n6759), .B(n6760), .C(n6761), .D(n6762), .Y(n6078) );
  AOI2BB2X1TS U6399 ( .B0(n11688), .B1(n6764), .A0N(n11361), .A1N(n5831), .Y(
        n6760) );
  NAND2X1TS U6401 ( .A(n10432), .B(n10428), .Y(n6764) );
  NAND4X1TS U6403 ( .A(n6077), .B(n5689), .C(n6765), .D(n6766), .Y(n6192) );
  NAND2X1TS U6422 ( .A(n11269), .B(n10994), .Y(n5490) );
  NAND2X1TS U6432 ( .A(n10162), .B(n10458), .Y(n5332) );
  NAND2X1TS U6433 ( .A(n12581), .B(n10995), .Y(n6450) );
  NAND2X1TS U6439 ( .A(n11264), .B(n11385), .Y(n5474) );
  NOR4XLTS U6444 ( .A(n6417), .B(n5878), .C(n5487), .D(n5833), .Y(n6091) );
  NAND2X1TS U6469 ( .A(n12217), .B(n10162), .Y(n6435) );
  NAND2X1TS U6472 ( .A(n11247), .B(n11409), .Y(n5877) );
  NAND2X1TS U6477 ( .A(n10884), .B(n12266), .Y(n6403) );
  NAND2X1TS U6511 ( .A(n9836), .B(n9326), .Y(n6779) );
  NAND2X1TS U6525 ( .A(sa12[4]), .B(n6793), .Y(n5701) );
  NAND2X1TS U6531 ( .A(n9443), .B(n9439), .Y(n5693) );
  NAND2X1TS U6538 ( .A(n10072), .B(n10075), .Y(n6792) );
  NAND2X1TS U6546 ( .A(n9431), .B(n9836), .Y(n6785) );
  NAND2X1TS U6553 ( .A(n12256), .B(n9961), .Y(n6503) );
  NOR4XLTS U6555 ( .A(n6806), .B(n6807), .C(n6808), .D(n6809), .Y(n5707) );
  NAND2X1TS U6557 ( .A(n10869), .B(n10913), .Y(n6474) );
  NAND2X1TS U6558 ( .A(n11710), .B(n12521), .Y(n6481) );
  NAND2X1TS U6582 ( .A(n10448), .B(n9774), .Y(n6498) );
  NAND4X1TS U6583 ( .A(n6817), .B(n6818), .C(n6819), .D(n6820), .Y(n6122) );
  AOI2BB2X1TS U6594 ( .B0(n11706), .B1(n6822), .A0N(n11367), .A1N(n5887), .Y(
        n6818) );
  NAND2X1TS U6596 ( .A(n10449), .B(n10445), .Y(n6822) );
  NAND4X1TS U6598 ( .A(n6121), .B(n5714), .C(n6823), .D(n6824), .Y(n6232) );
  NAND2X1TS U6617 ( .A(n11317), .B(n11006), .Y(n5556) );
  NAND2X1TS U6627 ( .A(n10170), .B(n10465), .Y(n5371) );
  NAND2X1TS U6628 ( .A(n12590), .B(n11007), .Y(n6522) );
  NAND2X1TS U6634 ( .A(n11312), .B(n11391), .Y(n5540) );
  NOR4XLTS U6639 ( .A(n6489), .B(n5934), .C(n5553), .D(n5889), .Y(n6135) );
  NAND2X1TS U6659 ( .A(n10542), .B(n10445), .Y(n6133) );
  NAND2X1TS U6664 ( .A(n12241), .B(n10169), .Y(n6507) );
  NAND2X1TS U6667 ( .A(n11295), .B(n11413), .Y(n5933) );
  NAND2X1TS U6672 ( .A(n10914), .B(n12274), .Y(n6475) );
  NAND2X1TS U6706 ( .A(n9880), .B(n9343), .Y(n6837) );
  NAND2X1TS U6720 ( .A(sa23[4]), .B(n6851), .Y(n5726) );
  NAND2X1TS U6726 ( .A(n9545), .B(n9541), .Y(n5718) );
  NAND2X1TS U6733 ( .A(n10100), .B(n10103), .Y(n6850) );
  NAND2X1TS U6741 ( .A(n9534), .B(n9880), .Y(n6843) );
  NOR4XLTS U6744 ( .A(n6860), .B(n6861), .C(n6862), .D(n6863), .Y(n6859) );
  NAND2X1TS U6755 ( .A(n11760), .B(n11331), .Y(n6616) );
  NOR4XLTS U6761 ( .A(n5758), .B(n6869), .C(n6870), .D(n6871), .Y(n5977) );
  NAND2X1TS U6767 ( .A(n11018), .B(n9711), .Y(n6372) );
  NAND4X1TS U6772 ( .A(n6876), .B(n6877), .C(n6878), .D(n6879), .Y(n6875) );
  NOR4XLTS U6773 ( .A(n5643), .B(n5978), .C(n5949), .D(n6880), .Y(n6879) );
  NAND2X1TS U6776 ( .A(n11758), .B(n10202), .Y(n6672) );
  NAND2X1TS U6777 ( .A(n6882), .B(n6883), .Y(n5949) );
  NAND2X1TS U6783 ( .A(n12062), .B(n10576), .Y(n6673) );
  NAND2X1TS U6785 ( .A(n10546), .B(n10577), .Y(n6620) );
  NAND2X1TS U6790 ( .A(n12054), .B(n11740), .Y(n6610) );
  NAND2X1TS U6795 ( .A(n12543), .B(n11758), .Y(n6630) );
  NAND2X1TS U6799 ( .A(n6334), .B(n12004), .Y(n5955) );
  NAND2X1TS U6801 ( .A(n10546), .B(n12279), .Y(n6664) );
  NOR4XLTS U6802 ( .A(n5766), .B(n5757), .C(n6894), .D(n6895), .Y(n6893) );
  NAND2X1TS U6804 ( .A(n10549), .B(n11353), .Y(n6364) );
  NAND2X1TS U6821 ( .A(n10233), .B(n10518), .Y(n6617) );
  AOI2BB2X1TS U6826 ( .B0(n10178), .B1(n6286), .A0N(n9781), .A1N(n6374), .Y(
        n6876) );
  OAI221XLTS U6832 ( .A0(n11736), .A1(n10197), .B0(n10518), .B1(n11746), .C0(
        n5963), .Y(n6874) );
  NAND2X1TS U6835 ( .A(n12544), .B(n10947), .Y(n6345) );
  NAND2X1TS U6838 ( .A(n10976), .B(n10518), .Y(n6295) );
  NAND2X1TS U6839 ( .A(n10230), .B(n11982), .Y(n6649) );
  NAND2X1TS U6857 ( .A(n6334), .B(n9778), .Y(n5586) );
  NAND2X1TS U6861 ( .A(n12681), .B(n6906), .Y(n5662) );
  NAND2X1TS U6863 ( .A(n11349), .B(n12537), .Y(n6340) );
  NAND3X1TS U6903 ( .A(n12681), .B(n6904), .C(n9344), .Y(n6277) );
  NAND2X1TS U6907 ( .A(sa01[4]), .B(n9345), .Y(n6637) );
  NAND2X1TS U6917 ( .A(n10048), .B(n6917), .Y(n6897) );
  NAND2X1TS U6919 ( .A(n10721), .B(n6918), .Y(n6338) );
  NAND2X1TS U6922 ( .A(n12680), .B(n6318), .Y(n6351) );
  NAND2X1TS U6925 ( .A(n5974), .B(n11329), .Y(n6648) );
  NAND2X1TS U6927 ( .A(sa01[6]), .B(n9824), .Y(n6317) );
  NAND2X1TS U6931 ( .A(n10229), .B(n10226), .Y(n5974) );
  NAND2X1TS U6934 ( .A(n10722), .B(sa01[5]), .Y(n6640) );
  NAND2X1TS U6935 ( .A(sa01[0]), .B(sa01[3]), .Y(n6872) );
  XNOR2X1TS U6941 ( .A(w2[31]), .B(n6919), .Y(N151) );
  OAI2BB2XLTS U6942 ( .B0(text_in_r[63]), .B1(n12696), .A0N(n6920), .A1N(
        n12717), .Y(n6919) );
  XNOR2X1TS U6946 ( .A(w2[30]), .B(n6928), .Y(N150) );
  OAI2BB2XLTS U6947 ( .B0(text_in_r[62]), .B1(n12697), .A0N(n6929), .A1N(
        n12715), .Y(n6928) );
  XNOR2X1TS U6951 ( .A(w2[29]), .B(n6937), .Y(N149) );
  OAI2BB2XLTS U6952 ( .B0(text_in_r[61]), .B1(n12698), .A0N(n6938), .A1N(
        n12719), .Y(n6937) );
  AOI2BB2X1TS U6953 ( .B0(n6939), .B1(n6940), .A0N(n6939), .A1N(n6940), .Y(
        n6938) );
  OAI2BB2XLTS U6957 ( .B0(text_in_r[60]), .B1(n9519), .A0N(n9518), .A1N(
        text_in_r[60]), .Y(n6945) );
  XOR2X1TS U6958 ( .A(n6946), .B(n6947), .Y(n6944) );
  XOR2X1TS U6959 ( .A(n6948), .B(n6949), .Y(n6947) );
  OAI2BB2XLTS U6965 ( .B0(text_in_r[59]), .B1(n9514), .A0N(n9513), .A1N(
        text_in_r[59]), .Y(n6955) );
  XOR2X1TS U6966 ( .A(n6956), .B(n6957), .Y(n6954) );
  XOR2X1TS U6967 ( .A(n6958), .B(n6959), .Y(n6957) );
  XNOR2X1TS U6974 ( .A(w2[26]), .B(n6961), .Y(N146) );
  OAI2BB2XLTS U6975 ( .B0(text_in_r[58]), .B1(n12700), .A0N(n6962), .A1N(
        n12714), .Y(n6961) );
  AOI2BB2X1TS U6976 ( .B0(n9783), .B1(n6963), .A0N(n9783), .A1N(n6963), .Y(
        n6962) );
  XNOR2X1TS U6977 ( .A(n1286), .B(n6964), .Y(n6963) );
  OAI2BB2XLTS U6980 ( .B0(text_in_r[57]), .B1(n9509), .A0N(n9508), .A1N(
        text_in_r[57]), .Y(n6967) );
  XOR2X1TS U6981 ( .A(n6968), .B(n6969), .Y(n6966) );
  XOR2X1TS U6982 ( .A(n6970), .B(n6971), .Y(n6969) );
  XNOR2X1TS U6988 ( .A(w2[24]), .B(n6973), .Y(N144) );
  OAI2BB2XLTS U6989 ( .B0(text_in_r[56]), .B1(n12701), .A0N(n6974), .A1N(
        n12718), .Y(n6973) );
  AOI2BB2X1TS U6990 ( .B0(n1303), .B1(n6975), .A0N(n1303), .A1N(n6975), .Y(
        n6974) );
  XNOR2X1TS U6992 ( .A(w2[23]), .B(n6977), .Y(N135) );
  OAI2BB2XLTS U6993 ( .B0(text_in_r[55]), .B1(n12702), .A0N(n6978), .A1N(
        n12715), .Y(n6977) );
  AOI2BB2X1TS U6994 ( .B0(n6934), .B1(n6979), .A0N(n6934), .A1N(n6979), .Y(
        n6978) );
  XNOR2X1TS U6997 ( .A(w2[22]), .B(n6981), .Y(N134) );
  OAI2BB2XLTS U6998 ( .B0(text_in_r[54]), .B1(n12703), .A0N(n6982), .A1N(
        n12714), .Y(n6981) );
  AOI2BB2X1TS U6999 ( .B0(n6941), .B1(n6983), .A0N(n6941), .A1N(n6983), .Y(
        n6982) );
  XNOR2X1TS U7002 ( .A(w2[21]), .B(n6987), .Y(N133) );
  OAI2BB2XLTS U7003 ( .B0(text_in_r[53]), .B1(n12703), .A0N(n6988), .A1N(
        n12714), .Y(n6987) );
  AOI2BB2X1TS U7004 ( .B0(n6951), .B1(n6989), .A0N(n6951), .A1N(n6989), .Y(
        n6988) );
  OAI2BB2XLTS U7007 ( .B0(text_in_r[52]), .B1(n9504), .A0N(n9503), .A1N(
        text_in_r[52]), .Y(n6993) );
  XOR2X1TS U7008 ( .A(n6994), .B(n6995), .Y(n6992) );
  XNOR2X1TS U7009 ( .A(n1278), .B(n6996), .Y(n6995) );
  OAI2BB2XLTS U7015 ( .B0(text_in_r[51]), .B1(n9499), .A0N(n9498), .A1N(
        text_in_r[51]), .Y(n7003) );
  XOR2X1TS U7016 ( .A(n7004), .B(n7005), .Y(n7002) );
  XNOR2X1TS U7017 ( .A(n7006), .B(n6999), .Y(n7005) );
  XNOR2X1TS U7023 ( .A(w2[18]), .B(n7010), .Y(N130) );
  OAI2BB2XLTS U7024 ( .B0(text_in_r[50]), .B1(n12705), .A0N(n7011), .A1N(
        n12716), .Y(n7010) );
  AOI2BB2X1TS U7025 ( .B0(n12662), .B1(n7012), .A0N(n1271), .A1N(n7012), .Y(
        n7011) );
  XNOR2X1TS U7026 ( .A(n9178), .B(n1297), .Y(n7012) );
  XNOR2X1TS U7028 ( .A(n1558), .B(n1598), .Y(n1298) );
  OAI2BB2XLTS U7030 ( .B0(text_in_r[49]), .B1(n9495), .A0N(n9494), .A1N(
        text_in_r[49]), .Y(n7014) );
  XOR2X1TS U7031 ( .A(n7015), .B(n7016), .Y(n7013) );
  XNOR2X1TS U7032 ( .A(n7017), .B(n6999), .Y(n7016) );
  XNOR2X1TS U7039 ( .A(w2[16]), .B(n7020), .Y(N128) );
  OAI2BB2XLTS U7040 ( .B0(text_in_r[48]), .B1(n12707), .A0N(n7021), .A1N(
        n12716), .Y(n7020) );
  AOI2BB2X1TS U7041 ( .B0(n12663), .B1(n7022), .A0N(n1292), .A1N(n7022), .Y(
        n7021) );
  XNOR2X1TS U7042 ( .A(n7019), .B(n7000), .Y(n7022) );
  XNOR2X1TS U7045 ( .A(w2[15]), .B(n7024), .Y(N119) );
  OAI2BB2XLTS U7046 ( .B0(text_in_r[47]), .B1(n12707), .A0N(n7025), .A1N(
        n12714), .Y(n7024) );
  AOI2BB2X1TS U7047 ( .B0(n7026), .B1(n7027), .A0N(n7026), .A1N(n7027), .Y(
        n7025) );
  XNOR2X1TS U7051 ( .A(w2[14]), .B(n7029), .Y(N118) );
  OAI2BB2XLTS U7052 ( .B0(text_in_r[46]), .B1(n12708), .A0N(n7030), .A1N(
        n12718), .Y(n7029) );
  AOI2BB2X1TS U7053 ( .B0(n7031), .B1(n7032), .A0N(n7031), .A1N(n7032), .Y(
        n7030) );
  XNOR2X1TS U7056 ( .A(w2[13]), .B(n7033), .Y(N117) );
  OAI2BB2XLTS U7057 ( .B0(text_in_r[45]), .B1(n12709), .A0N(n7034), .A1N(
        n12715), .Y(n7033) );
  AOI2BB2X1TS U7058 ( .B0(n9459), .B1(n7035), .A0N(n9460), .A1N(n7035), .Y(
        n7034) );
  XNOR2X1TS U7059 ( .A(n6997), .B(n7036), .Y(n7035) );
  OAI2BB2XLTS U7062 ( .B0(text_in_r[44]), .B1(n9489), .A0N(n9489), .A1N(
        text_in_r[44]), .Y(n7038) );
  XOR2X1TS U7063 ( .A(n7039), .B(n7040), .Y(n7037) );
  XOR2X1TS U7064 ( .A(n7041), .B(n7042), .Y(n7040) );
  XNOR2X1TS U7067 ( .A(n1562), .B(n9490), .Y(n7039) );
  NAND4BX1TS U7070 ( .AN(n7047), .B(n7048), .C(n7049), .D(n7050), .Y(n7046) );
  OAI222X1TS U7078 ( .A0(n11778), .A1(n8135), .B0(n12070), .B1(n10601), .C0(
        n7080), .C1(n11438), .Y(n7047) );
  NAND4BX1TS U7079 ( .AN(n7082), .B(n7083), .C(n7084), .D(n7085), .Y(n7045) );
  OAI2BB2XLTS U7083 ( .B0(text_in_r[43]), .B1(n9485), .A0N(n9484), .A1N(
        text_in_r[43]), .Y(n7093) );
  XOR2X1TS U7084 ( .A(n7094), .B(n7095), .Y(n7092) );
  XNOR2X1TS U7085 ( .A(n7096), .B(n1604), .Y(n7095) );
  NAND4BX1TS U7088 ( .AN(n7101), .B(n7102), .C(n7103), .D(n7104), .Y(n7100) );
  OAI222X1TS U7096 ( .A0(n12094), .A1(n8069), .B0(n12304), .B1(n11043), .C0(
        n7134), .C1(n11808), .Y(n7101) );
  NAND4BX1TS U7097 ( .AN(n7136), .B(n7137), .C(n7138), .D(n7139), .Y(n7099) );
  XNOR2X1TS U7102 ( .A(n9177), .B(n7146), .Y(n7094) );
  OAI222X1TS U7113 ( .A0(n11468), .A1(n11832), .B0(n11838), .B1(n11427), .C0(
        n10618), .C1(n10010), .Y(n7168) );
  XNOR2X1TS U7122 ( .A(w2[10]), .B(n7192), .Y(N114) );
  OAI2BB2XLTS U7123 ( .B0(text_in_r[42]), .B1(n12707), .A0N(n7193), .A1N(
        n12715), .Y(n7192) );
  XNOR2X1TS U7125 ( .A(n1601), .B(n7195), .Y(n7194) );
  NAND3X1TS U7127 ( .A(n7196), .B(n7197), .C(n7198), .Y(n1560) );
  NOR4XLTS U7128 ( .A(n7199), .B(n7200), .C(n7201), .D(n7202), .Y(n7197) );
  NOR4XLTS U7132 ( .A(n7210), .B(n7211), .C(n7212), .D(n7213), .Y(n7196) );
  AO22X1TS U7133 ( .A0(n7214), .A1(n12455), .B0(n11432), .B1(n7215), .Y(n7213)
         );
  NAND4X1TS U7138 ( .A(n7223), .B(n7138), .C(n7224), .D(n7225), .Y(n7222) );
  XNOR2X1TS U7153 ( .A(n9220), .B(n1284), .Y(n1271) );
  OAI2BB2XLTS U7176 ( .B0(text_in_r[41]), .B1(n9480), .A0N(n9479), .A1N(
        text_in_r[41]), .Y(n7341) );
  XOR2X1TS U7177 ( .A(n7342), .B(n7343), .Y(n7340) );
  XOR2X1TS U7178 ( .A(n7344), .B(n7345), .Y(n7343) );
  NAND3X1TS U7181 ( .A(n7346), .B(n7347), .C(n7348), .Y(n1600) );
  NOR4XLTS U7182 ( .A(n7349), .B(n7350), .C(n7351), .D(n7352), .Y(n7348) );
  NOR4XLTS U7186 ( .A(n7360), .B(n7361), .C(n7362), .D(n7363), .Y(n7347) );
  NOR4XLTS U7192 ( .A(n7373), .B(n7374), .C(n7375), .D(n7376), .Y(n7372) );
  AOI2BB2X1TS U7200 ( .B0(n11055), .B1(n7395), .A0N(n7180), .A1N(n11796), .Y(
        n7386) );
  OAI33XLTS U7205 ( .A0(n8666), .A1(n11842), .A2(n7404), .B0(n9496), .B1(
        n10298), .B2(sa20[4]), .Y(n7399) );
  NAND2X1TS U7207 ( .A(n12109), .B(n11547), .Y(n7206) );
  NAND3X1TS U7241 ( .A(n7470), .B(n7471), .C(n7472), .Y(n1513) );
  NOR4XLTS U7243 ( .A(n7477), .B(n7478), .C(n7479), .D(n7480), .Y(n7471) );
  XNOR2X1TS U7249 ( .A(w2[8]), .B(n7498), .Y(N112) );
  OAI2BB2XLTS U7250 ( .B0(text_in_r[40]), .B1(n12712), .A0N(n7499), .A1N(
        n12716), .Y(n7498) );
  AOI2BB2X1TS U7251 ( .B0(n1292), .B1(n7500), .A0N(n1292), .A1N(n7500), .Y(
        n7499) );
  XNOR2X1TS U7252 ( .A(n6972), .B(n9793), .Y(n7500) );
  XNOR2X1TS U7254 ( .A(n1568), .B(n7028), .Y(n6926) );
  NAND4X1TS U7259 ( .A(n7506), .B(n7137), .C(n7507), .D(n7508), .Y(n7505) );
  NOR4XLTS U7275 ( .A(n7353), .B(n7540), .C(n7541), .D(n7542), .Y(n7112) );
  OAI33XLTS U7278 ( .A0(n9842), .A1(n12322), .A2(n7547), .B0(n9841), .B1(
        n11128), .B2(sa13[4]), .Y(n7541) );
  NAND2X1TS U7288 ( .A(n10025), .B(n10688), .Y(n7370) );
  XNOR2X1TS U7292 ( .A(n6976), .B(n9779), .Y(n1292) );
  NAND4X1TS U7301 ( .A(n7595), .B(n7596), .C(n7597), .D(n7598), .Y(n7264) );
  NAND4X1TS U7303 ( .A(n7602), .B(n7603), .C(n7604), .D(n7605), .Y(n7601) );
  AND4X1TS U7310 ( .A(n7615), .B(n7616), .C(n7617), .D(n7618), .Y(n7597) );
  NOR4XLTS U7319 ( .A(n7636), .B(n7637), .C(n7638), .D(n7639), .Y(n7635) );
  NAND4X1TS U7320 ( .A(n7640), .B(n7641), .C(n7642), .D(n7643), .Y(n7639) );
  AO22X1TS U7329 ( .A0(n7330), .A1(n12618), .B0(n7665), .B1(n11591), .Y(n7637)
         );
  XNOR2X1TS U7342 ( .A(w2[7]), .B(n7701), .Y(N103) );
  OAI2BB2XLTS U7343 ( .B0(text_in_r[39]), .B1(n12712), .A0N(n7702), .A1N(
        n12717), .Y(n7701) );
  XNOR2X1TS U7345 ( .A(n6953), .B(n6985), .Y(n7703) );
  NAND4X1TS U7350 ( .A(n7483), .B(n7708), .C(n7709), .D(n7710), .Y(n7707) );
  OA22X1TS U7355 ( .A0(n10660), .A1(n9861), .B0(n12356), .B1(n7496), .Y(n7714)
         );
  NOR4XLTS U7357 ( .A(n7717), .B(n7718), .C(n7719), .D(n7720), .Y(n7483) );
  NAND3X1TS U7358 ( .A(n7721), .B(n7722), .C(n7723), .Y(n7720) );
  OA22X1TS U7361 ( .A0(n9520), .A1(n11868), .B0(n7729), .B1(n12357), .Y(n7721)
         );
  XNOR2X1TS U7372 ( .A(n9127), .B(n9151), .Y(n6953) );
  NAND2X1TS U7378 ( .A(n11474), .B(n12089), .Y(n7561) );
  NAND2X1TS U7381 ( .A(n11568), .B(n10320), .Y(n7104) );
  NOR4XLTS U7386 ( .A(n7758), .B(n7759), .C(n7760), .D(n7761), .Y(n7354) );
  NOR4XLTS U7399 ( .A(n7423), .B(n7780), .C(n7781), .D(n7782), .Y(n7779) );
  NAND2X1TS U7401 ( .A(n12109), .B(n9801), .Y(n7380) );
  NAND2X1TS U7404 ( .A(n11878), .B(n10673), .Y(n7050) );
  NAND2X1TS U7408 ( .A(n11541), .B(n10038), .Y(n7788) );
  NOR4XLTS U7409 ( .A(n7790), .B(n7791), .C(n7792), .D(n7793), .Y(n7203) );
  XNOR2X1TS U7420 ( .A(w2[6]), .B(n7805), .Y(N102) );
  OAI2BB2XLTS U7421 ( .B0(text_in_r[38]), .B1(n12712), .A0N(n7806), .A1N(
        n12718), .Y(n7805) );
  XNOR2X1TS U7423 ( .A(n6936), .B(n9460), .Y(n7807) );
  NAND4X1TS U7430 ( .A(n7817), .B(n7818), .C(n7819), .D(n7820), .Y(n7633) );
  NOR4XLTS U7437 ( .A(n7478), .B(n7830), .C(n7831), .D(n7832), .Y(n7808) );
  OAI2BB2XLTS U7439 ( .B0(n7835), .B1(n7739), .A0N(n7836), .A1N(n11151), .Y(
        n7831) );
  OAI2BB2XLTS U7440 ( .B0(n11529), .B1(n7837), .A0N(n11926), .A1N(n7838), .Y(
        n7830) );
  AO22X1TS U7441 ( .A0(n11156), .A1(n12143), .B0(n9542), .B1(n7682), .Y(n7478)
         );
  OAI33XLTS U7453 ( .A0(n11523), .A1(n9873), .A2(n7860), .B0(n9374), .B1(n9874), .B2(n11904), .Y(n7852) );
  OAI222X1TS U7454 ( .A0(n10065), .A1(n10338), .B0(n11598), .B1(n10646), .C0(
        n11558), .C1(n10724), .Y(n7851) );
  NAND2X1TS U7469 ( .A(n10022), .B(n9818), .Y(n7128) );
  NAND4X1TS U7472 ( .A(n7874), .B(n7875), .C(n7876), .D(n7877), .Y(n7350) );
  NAND2X1TS U7475 ( .A(n10623), .B(n11076), .Y(n7531) );
  NAND2X1TS U7479 ( .A(n9471), .B(n10257), .Y(n7563) );
  NAND4X1TS U7481 ( .A(n7883), .B(n7884), .C(n7885), .D(n7886), .Y(n7742) );
  NOR4XLTS U7482 ( .A(n7349), .B(n7887), .C(n7888), .D(n7889), .Y(n7886) );
  NAND4BX1TS U7487 ( .AN(n7894), .B(n7895), .C(n7896), .D(n7897), .Y(n7349) );
  NOR4XLTS U7488 ( .A(n7898), .B(n7899), .C(n7900), .D(n7901), .Y(n7896) );
  NAND2X1TS U7496 ( .A(n12321), .B(n11043), .Y(n7564) );
  NAND2X1TS U7499 ( .A(n10328), .B(n12462), .Y(n7765) );
  NOR4XLTS U7503 ( .A(n7911), .B(n7912), .C(n7913), .D(n7914), .Y(n7910) );
  NAND2X1TS U7512 ( .A(n9467), .B(n10009), .Y(n7074) );
  NAND4X1TS U7515 ( .A(n7921), .B(n7922), .C(n7923), .D(n7924), .Y(n7200) );
  NAND2X1TS U7518 ( .A(n11049), .B(n10614), .Y(n7421) );
  NAND2X1TS U7522 ( .A(n10013), .B(n12629), .Y(n7385) );
  NAND4X1TS U7524 ( .A(n7930), .B(n7931), .C(n7932), .D(n7933), .Y(n7773) );
  NOR4XLTS U7525 ( .A(n7199), .B(n7934), .C(n7935), .D(n7936), .Y(n7933) );
  NAND4BX1TS U7530 ( .AN(n7941), .B(n7942), .C(n7943), .D(n7944), .Y(n7199) );
  NOR4XLTS U7531 ( .A(n7945), .B(n7946), .C(n7947), .D(n7948), .Y(n7943) );
  NAND2X1TS U7539 ( .A(n11843), .B(n10601), .Y(n7395) );
  NAND2X1TS U7542 ( .A(n10037), .B(n11770), .Y(n7797) );
  NAND2X1TS U7553 ( .A(n10089), .B(n10691), .Y(n7289) );
  XNOR2X1TS U7563 ( .A(w2[5]), .B(n7994), .Y(N101) );
  OAI2BB2XLTS U7564 ( .B0(text_in_r[37]), .B1(n12712), .A0N(n7995), .A1N(
        n12719), .Y(n7994) );
  XNOR2X1TS U7566 ( .A(n6942), .B(n6998), .Y(n7996) );
  XNOR2X1TS U7568 ( .A(n1519), .B(n1643), .Y(n7001) );
  NAND4X1TS U7571 ( .A(n7708), .B(n8000), .C(n8001), .D(n8002), .Y(n7999) );
  NAND2X1TS U7576 ( .A(n11523), .B(n10723), .Y(n7664) );
  NAND4X1TS U7579 ( .A(n8007), .B(n8008), .C(n8009), .D(n8010), .Y(n8006) );
  AOI2BB2X1TS U7587 ( .B0(n12618), .B1(n7665), .A0N(n10646), .A1N(n7494), .Y(
        n8011) );
  NAND4X1TS U7588 ( .A(n8015), .B(n8016), .C(n8017), .D(n8018), .Y(n7477) );
  NOR4XLTS U7589 ( .A(n8019), .B(n8020), .C(n7704), .D(n8021), .Y(n8018) );
  NAND2X1TS U7591 ( .A(n9866), .B(n10282), .Y(n7643) );
  NAND4X1TS U7592 ( .A(n8023), .B(n8024), .C(n8025), .D(n8026), .Y(n7704) );
  NOR4XLTS U7599 ( .A(n7311), .B(n7857), .C(n8029), .D(n8030), .Y(n8017) );
  NOR4XLTS U7624 ( .A(n8051), .B(n8052), .C(n8053), .D(n8054), .Y(n7562) );
  NOR4XLTS U7630 ( .A(n8058), .B(n7360), .C(n8059), .D(n8060), .Y(n8038) );
  OAI2BB2XLTS U7638 ( .B0(n7125), .B1(n11932), .A0N(n8065), .A1N(n7526), .Y(
        n8064) );
  NAND4X1TS U7640 ( .A(n8066), .B(n8067), .C(n8068), .D(n7897), .Y(n7228) );
  NAND2X1TS U7641 ( .A(n10688), .B(n12088), .Y(n7897) );
  NAND2X1TS U7644 ( .A(n11533), .B(n10325), .Y(n7870) );
  NAND2X1TS U7645 ( .A(n11456), .B(n10025), .Y(n7877) );
  NAND4X1TS U7652 ( .A(n7502), .B(n8072), .C(n8073), .D(n8074), .Y(n7097) );
  NOR4XLTS U7653 ( .A(n7220), .B(n7511), .C(n8075), .D(n8076), .Y(n8074) );
  NAND4X1TS U7659 ( .A(n8079), .B(n8080), .C(n7356), .D(n8081), .Y(n7511) );
  NAND2X1TS U7660 ( .A(n10605), .B(n12312), .Y(n7356) );
  NAND2X1TS U7663 ( .A(n10605), .B(n10253), .Y(n7754) );
  NAND2X1TS U7664 ( .A(n12640), .B(n11078), .Y(n7768) );
  NAND4X1TS U7668 ( .A(n8086), .B(n8087), .C(n8088), .D(n7769), .Y(n7220) );
  NAND2X1TS U7669 ( .A(n10735), .B(n11473), .Y(n7769) );
  AOI222XLTS U7671 ( .A0(n11113), .A1(n12320), .B0(n11112), .B1(n11808), .C0(
        n12322), .C1(n12082), .Y(n8090) );
  NAND4X1TS U7687 ( .A(n8098), .B(n8099), .C(n8100), .D(n8101), .Y(n8097) );
  AOI2BB2X1TS U7690 ( .B0(n7253), .B1(n7878), .A0N(n12077), .A1N(n9830), .Y(
        n8099) );
  NAND2X1TS U7691 ( .A(n11933), .B(n11485), .Y(n7878) );
  NOR4XLTS U7708 ( .A(n8117), .B(n8118), .C(n8119), .D(n8120), .Y(n7379) );
  NOR4XLTS U7714 ( .A(n8124), .B(n7210), .C(n8125), .D(n8126), .Y(n8104) );
  OAI2BB2XLTS U7722 ( .B0(n7071), .B1(n11605), .A0N(n8131), .A1N(n12552), .Y(
        n8130) );
  NAND4X1TS U7724 ( .A(n8132), .B(n8133), .C(n8134), .D(n7944), .Y(n7156) );
  NAND2X1TS U7725 ( .A(n10670), .B(n12456), .Y(n7944) );
  NAND2X1TS U7728 ( .A(n7418), .B(n11547), .Y(n7916) );
  NAND2X1TS U7729 ( .A(n11788), .B(n11060), .Y(n7924) );
  NAND4X1TS U7736 ( .A(n7371), .B(n8138), .C(n8139), .D(n8140), .Y(n7043) );
  NOR4XLTS U7737 ( .A(n7148), .B(n7409), .C(n8141), .D(n8142), .Y(n8140) );
  NAND4X1TS U7744 ( .A(n8145), .B(n8146), .C(n7205), .D(n8147), .Y(n7409) );
  NAND2X1TS U7745 ( .A(n11025), .B(n12552), .Y(n7205) );
  NAND4X1TS U7747 ( .A(n8150), .B(n8151), .C(n7800), .D(n7785), .Y(n8149) );
  NAND2X1TS U7748 ( .A(n11027), .B(n10591), .Y(n7785) );
  NAND2X1TS U7749 ( .A(n11814), .B(n10614), .Y(n7800) );
  NAND4X1TS U7753 ( .A(n8152), .B(n8153), .C(n8154), .D(n7801), .Y(n7148) );
  NAND2X1TS U7754 ( .A(n11623), .B(n12109), .Y(n7801) );
  AOI222XLTS U7756 ( .A0(n11072), .A1(n11844), .B0(n11071), .B1(n11438), .C0(
        n11843), .C1(n11426), .Y(n8156) );
  NAND4X1TS U7772 ( .A(n8164), .B(n8165), .C(n8166), .D(n8167), .Y(n8163) );
  NAND2X1TS U7776 ( .A(n11603), .B(n11469), .Y(n7925) );
  NAND2X1TS U7785 ( .A(n10306), .B(n10642), .Y(n7978) );
  NAND4X1TS U7807 ( .A(n8212), .B(n8213), .C(n8214), .D(n8215), .Y(n7575) );
  OAI2BB2XLTS U7815 ( .B0(text_in_r[36]), .B1(n9475), .A0N(n9474), .A1N(
        text_in_r[36]), .Y(n8222) );
  XOR2X1TS U7817 ( .A(n8223), .B(n8224), .Y(n8221) );
  XNOR2X1TS U7818 ( .A(n7007), .B(n8225), .Y(n8224) );
  NAND2X1TS U7824 ( .A(n11945), .B(n10639), .Y(n7631) );
  NAND4X1TS U7843 ( .A(n8253), .B(n8254), .C(n8255), .D(n8256), .Y(n8252) );
  NAND4X1TS U7848 ( .A(n8257), .B(n8258), .C(n8259), .D(n7612), .Y(n8243) );
  NAND2X1TS U7851 ( .A(n11575), .B(n11652), .Y(n7593) );
  NAND2X1TS U7858 ( .A(n11183), .B(n10357), .Y(n7460) );
  NAND4X1TS U7859 ( .A(n8265), .B(n8266), .C(n8267), .D(n8201), .Y(n7955) );
  NAND2X1TS U7860 ( .A(n11134), .B(n11908), .Y(n8201) );
  OA22X1TS U7865 ( .A0(n12156), .A1(n10346), .B0(n8206), .B1(n11950), .Y(n8265) );
  XNOR2X1TS U7866 ( .A(n1275), .B(n1516), .Y(n7007) );
  NAND2X1TS U7874 ( .A(n8281), .B(n8282), .Y(n7669) );
  NAND2X1TS U7881 ( .A(n12183), .B(n7485), .Y(n8034) );
  NAND2X1TS U7893 ( .A(n10728), .B(n11593), .Y(n7482) );
  OAI2BB2XLTS U7895 ( .B0(n7659), .B1(n11598), .A0N(n9870), .A1N(n8296), .Y(
        n8295) );
  NAND4X1TS U7908 ( .A(n7301), .B(n7634), .C(n8307), .D(n8308), .Y(n7811) );
  NOR4XLTS U7909 ( .A(n7679), .B(n8309), .C(n8310), .D(n8311), .Y(n8308) );
  NOR4XLTS U7915 ( .A(n8316), .B(n8317), .C(n8318), .D(n8319), .Y(n8315) );
  NAND2X1TS U7922 ( .A(n9520), .B(n11510), .Y(n8286) );
  NAND4X1TS U7933 ( .A(n8330), .B(n8331), .C(n8332), .D(n8333), .Y(n8329) );
  NAND2X1TS U7935 ( .A(n12355), .B(n11922), .Y(n7665) );
  NAND2X1TS U7937 ( .A(n11902), .B(n10717), .Y(n7825) );
  NAND4X1TS U7941 ( .A(n8336), .B(n8337), .C(n8338), .D(n8339), .Y(n8335) );
  NAND2X1TS U7944 ( .A(n11102), .B(n10718), .Y(n8296) );
  NAND2X1TS U7948 ( .A(n9862), .B(n11529), .Y(n7838) );
  NAND2X1TS U7957 ( .A(n7986), .B(n11499), .Y(n7463) );
  AO22X1TS U7959 ( .A0(n12343), .A1(n7582), .B0(n10739), .B1(n8354), .Y(n8353)
         );
  NAND2X1TS U7965 ( .A(n10332), .B(n9516), .Y(n8259) );
  NAND2X1TS U7969 ( .A(n10701), .B(n11498), .Y(n7993) );
  NAND4X1TS U7990 ( .A(n7268), .B(n7578), .C(n7595), .D(n8379), .Y(n8168) );
  NOR4XLTS U8006 ( .A(n8390), .B(n8391), .C(n8392), .D(n8393), .Y(n7595) );
  NAND2X1TS U8009 ( .A(n9878), .B(n10086), .Y(n7296) );
  NAND2X1TS U8011 ( .A(n11087), .B(n11910), .Y(n8256) );
  NAND2X1TS U8018 ( .A(n11182), .B(n11188), .Y(n8216) );
  OAI2BB2XLTS U8020 ( .B0(n11165), .B1(n8270), .A0N(n7594), .A1N(n12636), .Y(
        n8401) );
  NAND2X1TS U8021 ( .A(n11199), .B(n12164), .Y(n7594) );
  NAND2X1TS U8028 ( .A(n10347), .B(n11119), .Y(n8240) );
  NAND2X1TS U8029 ( .A(n11187), .B(n11952), .Y(n8354) );
  NAND2X1TS U8039 ( .A(n10069), .B(n9869), .Y(n8305) );
  NAND4X1TS U8046 ( .A(n8426), .B(n8427), .C(n8428), .D(n8429), .Y(n7705) );
  NOR4XLTS U8047 ( .A(n7997), .B(n8029), .C(n7479), .D(n8430), .Y(n8429) );
  NAND4BX1TS U8048 ( .AN(n8322), .B(n8431), .C(n8432), .D(n8433), .Y(n8430) );
  NAND4X1TS U8053 ( .A(n8434), .B(n8435), .C(n8339), .D(n7855), .Y(n7479) );
  NAND2X1TS U8054 ( .A(n11854), .B(n9870), .Y(n7855) );
  NAND2X1TS U8055 ( .A(n11854), .B(n12487), .Y(n8339) );
  NAND2X1TS U8059 ( .A(n10082), .B(n12350), .Y(n8285) );
  OAI221XLTS U8060 ( .A0(n11107), .A1(n10286), .B0(n11559), .B1(n10073), .C0(
        n7848), .Y(n8436) );
  NAND2X1TS U8061 ( .A(n12632), .B(n11551), .Y(n7848) );
  NAND2X1TS U8064 ( .A(n11915), .B(n11956), .Y(n7684) );
  NAND2X1TS U8067 ( .A(n10728), .B(n12486), .Y(n8280) );
  NAND4X1TS U8071 ( .A(n8445), .B(n8446), .C(n8447), .D(n7328), .Y(n7997) );
  NAND2X1TS U8072 ( .A(n11156), .B(n11897), .Y(n7328) );
  NAND2X1TS U8086 ( .A(n11558), .B(n11107), .Y(n7491) );
  NAND2X1TS U8088 ( .A(n10062), .B(n9857), .Y(n8326) );
  NAND2X1TS U8095 ( .A(n9520), .B(n10337), .Y(n8340) );
  NOR4XLTS U8096 ( .A(n8020), .B(n7492), .C(n8455), .D(n8456), .Y(n8418) );
  NAND4X1TS U8101 ( .A(n8457), .B(n8458), .C(n8459), .D(n8460), .Y(n7492) );
  NAND2X1TS U8104 ( .A(n11956), .B(n11155), .Y(n8321) );
  NAND2X1TS U8105 ( .A(n10082), .B(n11898), .Y(n7845) );
  OAI2BB2XLTS U8109 ( .B0(n7690), .B1(n10652), .A0N(n12351), .A1N(n7663), .Y(
        n8461) );
  NAND2X1TS U8118 ( .A(n11867), .B(n11609), .Y(n7712) );
  NAND4X1TS U8122 ( .A(n8464), .B(n8465), .C(n8333), .D(n7849), .Y(n8020) );
  NAND2X1TS U8123 ( .A(n7682), .B(n12364), .Y(n7849) );
  NAND2X1TS U8125 ( .A(n12351), .B(n11861), .Y(n8333) );
  NAND2X1TS U8131 ( .A(n9552), .B(n10712), .Y(n7686) );
  NAND2X1TS U8142 ( .A(n10335), .B(n8470), .Y(n7829) );
  NAND4X1TS U8148 ( .A(n8471), .B(n8472), .C(n8473), .D(n8313), .Y(n8014) );
  NAND2X1TS U8149 ( .A(n11155), .B(n11592), .Y(n8313) );
  NAND2X1TS U8155 ( .A(n7847), .B(n11552), .Y(n7813) );
  NAND2X1TS U8164 ( .A(n10070), .B(n11151), .Y(n8284) );
  NAND2X1TS U8168 ( .A(n11860), .B(n11927), .Y(n7823) );
  NAND2X1TS U8191 ( .A(n10646), .B(n10711), .Y(n7332) );
  NAND2X1TS U8197 ( .A(sa31[0]), .B(n9370), .Y(n8466) );
  NAND2X1TS U8201 ( .A(n10341), .B(n9365), .Y(n7731) );
  NOR2BX1TS U8203 ( .AN(n9597), .B(n7730), .Y(n7836) );
  NAND2X1TS U8215 ( .A(n9366), .B(n10341), .Y(n8478) );
  NAND4X1TS U8231 ( .A(n8245), .B(n8483), .C(n8484), .D(n8485), .Y(n8482) );
  AOI2BB2X1TS U8239 ( .B0(n11093), .B1(n8490), .A0N(n11652), .A1N(n8491), .Y(
        n8261) );
  AOI2BB1X1TS U8242 ( .A0N(n7275), .A1N(n11188), .B0(n8386), .Y(n8493) );
  NAND2X1TS U8247 ( .A(n7446), .B(n10740), .Y(n8358) );
  NAND4X1TS U8249 ( .A(n8496), .B(n8497), .C(n8498), .D(n8373), .Y(n8494) );
  NAND2X1TS U8250 ( .A(n12637), .B(n12134), .Y(n8373) );
  NAND2X1TS U8251 ( .A(n11581), .B(n11172), .Y(n8498) );
  OAI221XLTS U8257 ( .A0(n11654), .A1(n11119), .B0(n11586), .B1(n10098), .C0(
        n8501), .Y(n8500) );
  NAND2X1TS U8260 ( .A(n10102), .B(n10739), .Y(n8398) );
  NAND2X1TS U8262 ( .A(n10697), .B(n11646), .Y(n7599) );
  NAND2X1TS U8265 ( .A(n10049), .B(n11640), .Y(n7451) );
  NAND2X1TS U8268 ( .A(n11505), .B(n12642), .Y(n8395) );
  NAND2X1TS U8273 ( .A(n10301), .B(n10701), .Y(n8189) );
  OA21XLTS U8290 ( .A0(n8521), .A1(n8522), .B0(n8400), .Y(n8518) );
  NAND2X1TS U8291 ( .A(n10101), .B(n11908), .Y(n8400) );
  NAND2X1TS U8295 ( .A(n11133), .B(n11193), .Y(n8363) );
  NAND2X1TS U8302 ( .A(n12165), .B(n10356), .Y(n7610) );
  NAND2X1TS U8304 ( .A(n11087), .B(n7467), .Y(n7574) );
  NAND2X1TS U8305 ( .A(n10750), .B(n11640), .Y(n7467) );
  NAND2X1TS U8313 ( .A(n12155), .B(n11653), .Y(n7979) );
  NAND2X1TS U8323 ( .A(n11641), .B(n9528), .Y(n8219) );
  NAND2X1TS U8326 ( .A(n11892), .B(n10050), .Y(n8385) );
  NAND2X1TS U8328 ( .A(n11493), .B(n10740), .Y(n8200) );
  NAND4X1TS U8332 ( .A(n8532), .B(n8533), .C(n8399), .D(n8188), .Y(n8531) );
  NAND2X1TS U8333 ( .A(n10101), .B(n12470), .Y(n8188) );
  NAND2X1TS U8335 ( .A(n12597), .B(n11091), .Y(n8399) );
  NAND4BX1TS U8351 ( .AN(n8396), .B(n8536), .C(n8537), .D(n8538), .Y(n8226) );
  NAND2X1TS U8358 ( .A(n10731), .B(n11174), .Y(n8521) );
  NAND2X1TS U8378 ( .A(n11180), .B(n10344), .Y(n8523) );
  NAND2X1TS U8386 ( .A(n9832), .B(n8546), .Y(n7454) );
  NAND2X1TS U8405 ( .A(n9832), .B(sa02[5]), .Y(n8488) );
  NAND2X1TS U8407 ( .A(n8525), .B(n8272), .Y(n8270) );
  NAND2X1TS U8409 ( .A(n9539), .B(n10731), .Y(n7630) );
  NAND2X1TS U8419 ( .A(n8525), .B(n9593), .Y(n8491) );
  XNOR2X1TS U8423 ( .A(n6997), .B(n1605), .Y(n6952) );
  NAND4BX1TS U8425 ( .AN(n7861), .B(n7746), .C(n7346), .D(n8547), .Y(n1607) );
  NOR4XLTS U8428 ( .A(n8551), .B(n8552), .C(n8553), .D(n8554), .Y(n7883) );
  AOI2BB2X1TS U8438 ( .B0(n11159), .B1(n7757), .A0N(n12113), .A1N(n7365), .Y(
        n8550) );
  NAND3X1TS U8439 ( .A(n8558), .B(n8559), .C(n8560), .Y(n8548) );
  OAI222X1TS U8442 ( .A0(n10266), .A1(n9838), .B0(n12319), .B1(n7229), .C0(
        n12464), .C1(n10022), .Y(n7556) );
  NAND2X1TS U8445 ( .A(n12119), .B(n12306), .Y(n7570) );
  NOR2BX1TS U8446 ( .AN(n10737), .B(n8562), .Y(n7757) );
  NAND4X1TS U8451 ( .A(n8565), .B(n8566), .C(n8567), .D(n8568), .Y(n8564) );
  NAND4X1TS U8453 ( .A(n8570), .B(n8571), .C(n8572), .D(n7544), .Y(n7887) );
  NAND2X1TS U8454 ( .A(n11569), .B(n11473), .Y(n7544) );
  NAND2X1TS U8465 ( .A(n11160), .B(n10057), .Y(n8043) );
  NAND2X1TS U8481 ( .A(n11038), .B(n10261), .Y(n8582) );
  NAND2X1TS U8485 ( .A(n10057), .B(n12314), .Y(n8056) );
  NAND2X1TS U8489 ( .A(n12639), .B(n11533), .Y(n8055) );
  NAND2X1TS U8492 ( .A(n11083), .B(n10686), .Y(n8080) );
  NAND2X1TS U8493 ( .A(n12319), .B(n11800), .Y(n7509) );
  NAND2X1TS U8502 ( .A(n10632), .B(n10257), .Y(n7567) );
  NAND2X1TS U8514 ( .A(n11534), .B(n11629), .Y(n8081) );
  NAND2X1TS U8521 ( .A(n10734), .B(n10686), .Y(n8063) );
  NAND2X1TS U8538 ( .A(n11535), .B(n7550), .Y(n7145) );
  NAND2X1TS U8542 ( .A(n10604), .B(n8047), .Y(n7256) );
  NOR4XLTS U8551 ( .A(n8607), .B(n8608), .C(n8609), .D(n8610), .Y(n8604) );
  NAND2X1TS U8563 ( .A(sa13[1]), .B(n11196), .Y(n8602) );
  NAND2X1TS U8567 ( .A(n11159), .B(n12090), .Y(n7236) );
  NAND2X1TS U8584 ( .A(n10738), .B(n9859), .Y(n8598) );
  NAND2X1TS U8593 ( .A(n9864), .B(n9867), .Y(n8578) );
  NAND2X1TS U8599 ( .A(n9860), .B(n10737), .Y(n8591) );
  NAND2X1TS U8601 ( .A(n10683), .B(n12307), .Y(n7523) );
  NAND2X1TS U8604 ( .A(n9868), .B(n9864), .Y(n8599) );
  NAND4BX1TS U8612 ( .AN(n7907), .B(n7777), .C(n7198), .D(n8614), .Y(n1565) );
  NOR4XLTS U8616 ( .A(n8618), .B(n8619), .C(n8620), .D(n8621), .Y(n7930) );
  NOR2BX1TS U8629 ( .AN(sa20[3]), .B(n8628), .Y(n7789) );
  AOI222XLTS U8632 ( .A0(n10269), .A1(n11621), .B0(n11938), .B1(n11546), .C0(
        n11066), .C1(n9801), .Y(n7381) );
  NAND4X1TS U8636 ( .A(n8632), .B(n8633), .C(n8634), .D(n8109), .Y(n8631) );
  NAND2X1TS U8637 ( .A(n11938), .B(n10290), .Y(n8109) );
  NAND4X1TS U8639 ( .A(n8636), .B(n8637), .C(n8638), .D(n7402), .Y(n7934) );
  NAND2X1TS U8640 ( .A(n11879), .B(n12107), .Y(n7402) );
  NAND2X1TS U8660 ( .A(n10289), .B(n12553), .Y(n8122) );
  NAND2X1TS U8666 ( .A(n11433), .B(n10002), .Y(n8646) );
  NAND2X1TS U8668 ( .A(n11765), .B(n11420), .Y(n8131) );
  NAND2X1TS U8679 ( .A(n11812), .B(n11066), .Y(n8121) );
  NAND2X1TS U8682 ( .A(n11461), .B(n10669), .Y(n8146) );
  NAND2X1TS U8688 ( .A(n11053), .B(n12630), .Y(n7389) );
  NAND2X1TS U8700 ( .A(n11065), .B(n11635), .Y(n8147) );
  NAND2X1TS U8707 ( .A(n11622), .B(n10668), .Y(n8129) );
  NAND2X1TS U8724 ( .A(n11066), .B(n11462), .Y(n7091) );
  NAND2X1TS U8728 ( .A(n11026), .B(n9575), .Y(n7184) );
  NOR4XLTS U8737 ( .A(n8672), .B(n8673), .C(n8674), .D(n8675), .Y(n8669) );
  NAND2X1TS U8753 ( .A(n11940), .B(n12456), .Y(n7164) );
  NAND2X1TS U8769 ( .A(n10705), .B(n9791), .Y(n8664) );
  NAND2X1TS U8779 ( .A(n10036), .B(n9795), .Y(n8679) );
  NAND2X1TS U8785 ( .A(n9792), .B(n10704), .Y(n8657) );
  NAND2X1TS U8787 ( .A(n10665), .B(n12070), .Y(n7435) );
  NAND2X1TS U8790 ( .A(n9796), .B(sa20[2]), .Y(n8665) );
  DFFQX1TS \sa13_reg[6]  ( .D(N70), .CK(clk), .Q(sa13[6]) );
  DFFQX1TS \sa13_reg[3]  ( .D(N67), .CK(clk), .Q(sa13[3]) );
  DFFQX1TS \sa02_reg[6]  ( .D(N150), .CK(clk), .Q(sa02[6]) );
  DFFQX1TS \sa01_reg[7]  ( .D(N215), .CK(clk), .Q(sa01[7]) );
  DFFQX1TS \sa33_reg[6]  ( .D(N38), .CK(clk), .Q(sa33[6]) );
  DFFQX1TS \sa10_reg[4]  ( .D(N260), .CK(clk), .Q(sa10[4]) );
  DFFQX1TS \sa21_reg[4]  ( .D(N180), .CK(clk), .Q(sa21[4]) );
  DFFQX1TS \sa30_reg[7]  ( .D(N231), .CK(clk), .Q(sa30[7]) );
  DFFQX1TS \sa00_reg[0]  ( .D(N272), .CK(clk), .Q(sa00[0]) );
  DFFQX1TS \sa33_reg[7]  ( .D(N39), .CK(clk), .Q(sa33[7]) );
  DFFQX1TS \sa23_reg[2]  ( .D(N50), .CK(clk), .Q(sa23[2]) );
  DFFQX1TS \sa22_reg[2]  ( .D(N114), .CK(clk), .Q(sa22[2]) );
  DFFQX1TS \sa12_reg[2]  ( .D(N130), .CK(clk), .Q(sa12[2]) );
  DFFQX1TS \sa11_reg[2]  ( .D(N194), .CK(clk), .Q(sa11[2]) );
  DFFQX1TS \sa33_reg[3]  ( .D(N35), .CK(clk), .Q(sa33[3]) );
  DFFQX1TS \sa30_reg[3]  ( .D(N227), .CK(clk), .Q(sa30[3]) );
  DFFQX1TS \sa20_reg[3]  ( .D(N243), .CK(clk), .Q(sa20[3]) );
  DFFQX1TS \sa02_reg[3]  ( .D(N147), .CK(clk), .Q(sa02[3]) );
  DFFQX1TS \sa02_reg[1]  ( .D(N145), .CK(clk), .Q(sa02[1]) );
  OAI32XLTS U4232 ( .A0(n10314), .A1(n9201), .A2(n12493), .B0(n4839), .B1(
        n10313), .Y(n4561) );
  OAI32XLTS U6112 ( .A0(n12680), .A1(n6637), .A2(n10230), .B0(n6638), .B1(
        n12680), .Y(n6365) );
  OAI32XLTS U2423 ( .A0(sa32[6]), .A1(n9045), .A2(n10955), .B0(n3099), .B1(
        n9852), .Y(n2615) );
  NOR2X1TS U8415 ( .A(n10344), .B(n11181), .Y(n8545) );
  AOI21X1TS U8031 ( .A0(n11890), .A1(n11576), .B0(n10045), .Y(n8406) );
  NOR2X1TS U8349 ( .A(n9877), .B(n12172), .Y(n8415) );
  NOR2X1TS U8279 ( .A(n11134), .B(n11491), .Y(n8413) );
  INVX2TS U8408 ( .A(n7630), .Y(n8272) );
  AOI211X1TS U8024 ( .A0(n12636), .A1(n8354), .B0(n8411), .C0(n8412), .Y(n8410) );
  OAI211X1TS U8023 ( .A0(n8408), .A1(n11586), .B0(n8409), .C0(n8410), .Y(n8407) );
  AOI211X1TS U8022 ( .A0(n10302), .A1(n10305), .B0(n8406), .C0(n8407), .Y(
        n7268) );
  NOR2X1TS U8361 ( .A(n10306), .B(n10639), .Y(n8175) );
  INVX2TS U8359 ( .A(n9565), .Y(n8364) );
  AOI22X1TS U8019 ( .A0(n11946), .A1(n11171), .B0(n11908), .B1(n12597), .Y(
        n8403) );
  INVX2TS U8404 ( .A(n8488), .Y(n8271) );
  NOR2X1TS U8016 ( .A(n11198), .B(n10745), .Y(n7973) );
  AOI211X1TS U8015 ( .A0(n11503), .A1(n8216), .B0(n8405), .C0(n7973), .Y(n8404) );
  OAI211X1TS U8014 ( .A0(n11187), .A1(n12171), .B0(n8403), .C0(n8404), .Y(
        n8402) );
  AOI211X1TS U8013 ( .A0(n10333), .A1(n9510), .B0(n8401), .C0(n8402), .Y(n7578) );
  NOR2X1TS U8248 ( .A(n11198), .B(n12170), .Y(n8390) );
  OAI211X1TS U8012 ( .A0(n11188), .A1(n10696), .B0(n8399), .C0(n8400), .Y(
        n8391) );
  NOR2X1TS U8411 ( .A(n10346), .B(n11640), .Y(n8396) );
  NOR2X1TS U8320 ( .A(n12156), .B(n11187), .Y(n8397) );
  AOI22X1TS U8004 ( .A0(n11944), .A1(n12478), .B0(n11497), .B1(n12595), .Y(
        n8389) );
  NOR2X1TS U8278 ( .A(n11133), .B(n12643), .Y(n8179) );
  AOI22X1TS U8000 ( .A0(n12596), .A1(n7300), .B0(n12471), .B1(n8370), .Y(n8382) );
  AOI22X1TS U7999 ( .A0(n11910), .A1(n12481), .B0(n10643), .B1(n9532), .Y(
        n8383) );
  NOR2X1TS U8243 ( .A(n11177), .B(n10357), .Y(n8386) );
  INVX2TS U7997 ( .A(n9482), .Y(n8190) );
  OAI22X1TS U7994 ( .A0(n8190), .A1(n11576), .B0(n7459), .B1(n11653), .Y(n8387) );
  AOI211X1TS U7991 ( .A0(n10332), .A1(n12642), .B0(n8380), .C0(n8381), .Y(
        n8379) );
  AOI22X1TS U7812 ( .A0(n10638), .A1(n12178), .B0(n12480), .B1(n9821), .Y(
        n8212) );
  AOI22X1TS U7811 ( .A0(n12177), .A1(n11172), .B0(n9629), .B1(n8187), .Y(n8213) );
  NOR2X1TS U8261 ( .A(n10045), .B(n11165), .Y(n8217) );
  AOI211X1TS U7808 ( .A0(n11909), .A1(n8216), .B0(n8217), .C0(n8218), .Y(n8215) );
  NOR2X1TS U7955 ( .A(n11193), .B(n12179), .Y(n8206) );
  NOR2X1TS U7989 ( .A(n11134), .B(n12479), .Y(n8250) );
  NOR2X1TS U7803 ( .A(n7465), .B(n10352), .Y(n7984) );
  NOR2X1TS U8355 ( .A(n12127), .B(n11639), .Y(n8204) );
  NOR2X1TS U7840 ( .A(n12162), .B(n11653), .Y(n8205) );
  AOI211X1TS U7802 ( .A0(n12136), .A1(n11946), .B0(n8204), .C0(n8205), .Y(
        n8195) );
  OAI211X1TS U7798 ( .A0(n12171), .A1(n11586), .B0(n8195), .C0(n8196), .Y(
        n8194) );
  AOI211X1TS U7797 ( .A0(n12643), .A1(n10739), .B0(n7984), .C0(n8194), .Y(
        n7596) );
  NOR2X1TS U7796 ( .A(n11892), .B(n7466), .Y(n7980) );
  NOR2X1TS U8299 ( .A(n11086), .B(n10639), .Y(n8182) );
  AOI22X1TS U7795 ( .A0(n11945), .A1(n7610), .B0(n10639), .B1(n9821), .Y(n8183) );
  OAI211X1TS U7791 ( .A0(n8182), .A1(n11178), .B0(n8183), .C0(n8184), .Y(n8181) );
  AOI211X1TS U7790 ( .A0(n12177), .A1(n12627), .B0(n7980), .C0(n8181), .Y(
        n7269) );
  AOI22X1TS U7789 ( .A0(n11908), .A1(n9532), .B0(n12641), .B1(n9822), .Y(n7457) );
  NOR2X1TS U7828 ( .A(n10346), .B(n10351), .Y(n8177) );
  NOR2X1TS U8796 ( .A(n10036), .B(n9795), .Y(n8648) );
  INVX2TS U8695 ( .A(n9561), .Y(n7404) );
  NOR2X1TS U8693 ( .A(n11788), .B(n11031), .Y(n8123) );
  NOR2X1TS U8756 ( .A(n9791), .B(n10705), .Y(n8667) );
  NOR2X1TS U8767 ( .A(n9799), .B(n9804), .Y(n8668) );
  NOR2X1TS U7779 ( .A(n10273), .B(n11432), .Y(n7065) );
  NOR2X1TS U7778 ( .A(n7065), .B(n10041), .Y(n7950) );
  NOR2X1TS U8783 ( .A(n9803), .B(n9800), .Y(n7154) );
  AOI22X1TS U7777 ( .A0(n11788), .A1(n11880), .B0(n11027), .B1(n11824), .Y(
        n8164) );
  NOR2X1TS U8658 ( .A(n11032), .B(n10269), .Y(n7786) );
  AOI22X1TS U7775 ( .A0(n11886), .A1(n7214), .B0(n11940), .B1(n7925), .Y(n8165) );
  AOI22X1TS U7773 ( .A0(n11824), .A1(n11462), .B0(n11622), .B1(n10674), .Y(
        n8167) );
  AOI22X1TS U7770 ( .A0(n11026), .A1(n11054), .B0(n9890), .B1(n11545), .Y(
        n8138) );
  NOR2X1TS U7768 ( .A(n11059), .B(n11782), .Y(n7802) );
  NOR2X1TS U7767 ( .A(n12107), .B(n10613), .Y(n7071) );
  INVX2TS U8786 ( .A(n7435), .Y(n7937) );
  OAI22X1TS U7765 ( .A0(n7937), .A1(n11468), .B0(n9813), .B1(n10599), .Y(n8161) );
  AOI211X1TS U7764 ( .A0(n9889), .A1(n7178), .B0(n8160), .C0(n8161), .Y(n8139)
         );
  NOR2X1TS U8634 ( .A(n10668), .B(n10014), .Y(n7069) );
  AOI22X1TS U7763 ( .A0(n11884), .A1(n8158), .B0(n7418), .B1(n12629), .Y(n8152) );
  NOR2X1TS U7762 ( .A(n11819), .B(n11438), .Y(n7945) );
  OAI22X1TS U7760 ( .A0(n11794), .A1(n11764), .B0(n11070), .B1(n11772), .Y(
        n8157) );
  AOI211X1TS U7759 ( .A0(n11061), .A1(n11066), .B0(n7945), .C0(n8157), .Y(
        n8153) );
  NOR2X1TS U7758 ( .A(n11790), .B(n10270), .Y(n7406) );
  AOI211X1TS U7755 ( .A0(n11825), .A1(n11633), .B0(n8155), .C0(n8156), .Y(
        n8154) );
  AOI211X1TS U7746 ( .A0(n11878), .A1(n11826), .B0(n8148), .C0(n8149), .Y(
        n8145) );
  AOI21X1TS U7743 ( .A0(n11766), .A1(n11771), .B0(n10664), .Y(n8141) );
  AOI22X1TS U7741 ( .A0(n10674), .A1(n12457), .B0(n11634), .B1(n12550), .Y(
        n8143) );
  AOI22X1TS U7739 ( .A0(n11623), .A1(n12551), .B0(n12631), .B1(n7067), .Y(
        n8144) );
  OAI211X1TS U7738 ( .A0(n11070), .A1(n10038), .B0(n8143), .C0(n8144), .Y(
        n8142) );
  AOI22X1TS U7735 ( .A0(n11824), .A1(n11060), .B0(n11031), .B1(n11431), .Y(
        n8132) );
  NOR2X1TS U7734 ( .A(n11938), .B(n10614), .Y(n7798) );
  NOR2X1TS U7731 ( .A(n11547), .B(n10290), .Y(n7180) );
  OAI22X1TS U7730 ( .A0(n9798), .A1(n10617), .B0(n7180), .B1(n11778), .Y(n8136) );
  OAI211X1TS U7727 ( .A0(n12329), .A1(n10294), .B0(n7924), .C0(n7916), .Y(
        n8137) );
  AOI211X1TS U7726 ( .A0(n11633), .A1(n11054), .B0(n8136), .C0(n8137), .Y(
        n8134) );
  NOR2X1TS U7723 ( .A(n10037), .B(n11439), .Y(n7941) );
  OAI211X1TS U7720 ( .A0(n12330), .A1(n11604), .B0(n8128), .C0(n8129), .Y(
        n8102) );
  OAI22X1TS U7718 ( .A0(n7937), .A1(n10595), .B0(n10664), .B1(n10599), .Y(
        n7210) );
  OAI22X1TS U7713 ( .A0(n11796), .A1(n10617), .B0(n10037), .B1(n11830), .Y(
        n8117) );
  OAI22X1TS U7712 ( .A0(n11778), .A1(n10293), .B0(n12148), .B1(n11772), .Y(
        n8118) );
  NOR2X1TS U8672 ( .A(n11783), .B(n12630), .Y(n7216) );
  NOR2X1TS U7710 ( .A(n11431), .B(n12455), .Y(n7425) );
  AOI22X1TS U7706 ( .A0(n11032), .A1(n10273), .B0(n10014), .B1(n7784), .Y(
        n8105) );
  NOR2X1TS U8625 ( .A(n11880), .B(n10290), .Y(n8110) );
  AOI22X1TS U7705 ( .A0(n11790), .A1(n11048), .B0(n11463), .B1(n10613), .Y(
        n8111) );
  NOR2X1TS U8758 ( .A(n10594), .B(n9463), .Y(n8114) );
  AOI211X1TS U7703 ( .A0(n9576), .A1(n11621), .B0(n8114), .C0(n8115), .Y(n8112) );
  OAI211X1TS U7702 ( .A0(n8110), .A1(n12330), .B0(n8111), .C0(n8112), .Y(n8106) );
  AOI22X1TS U7701 ( .A0(n11032), .A1(n11784), .B0(n11433), .B1(n10673), .Y(
        n8108) );
  OAI211X1TS U7700 ( .A0(n12327), .A1(n10595), .B0(n8108), .C0(n8109), .Y(
        n8107) );
  NOR2X1TS U7699 ( .A(n8106), .B(n8107), .Y(n7413) );
  INVX2TS U8562 ( .A(n8602), .Y(n8574) );
  NOR2X1TS U8609 ( .A(sa13[2]), .B(n9867), .Y(n8579) );
  NOR2X1TS U8607 ( .A(n11197), .B(n7528), .Y(n8590) );
  NOR2X1TS U8507 ( .A(n11455), .B(n11444), .Y(n8057) );
  NOR2X1TS U8570 ( .A(n9859), .B(n10737), .Y(n8600) );
  NOR2X1TS U8582 ( .A(n9871), .B(n9876), .Y(n8601) );
  NOR2X1TS U7694 ( .A(n10278), .B(n11038), .Y(n7119) );
  INVX2TS U8541 ( .A(n9556), .Y(n7547) );
  NOR2X1TS U7693 ( .A(n7119), .B(n9837), .Y(n7903) );
  NOR2X1TS U8597 ( .A(n9875), .B(n9872), .Y(n7226) );
  INVX2TS U8577 ( .A(n9841), .Y(n8603) );
  AOI22X1TS U7692 ( .A0(n11457), .A1(n11570), .B0(n10604), .B1(n11479), .Y(
        n8098) );
  OAI21X1TS U7689 ( .A0(n12640), .A1(n11628), .B0(n9886), .Y(n8100) );
  AOI22X1TS U7688 ( .A0(n11480), .A1(n11083), .B0(n10734), .B1(n10321), .Y(
        n8101) );
  AOI211X1TS U7686 ( .A0(n12638), .A1(n8096), .B0(n7903), .C0(n8097), .Y(n7502) );
  AOI22X1TS U7685 ( .A0(n7767), .A1(n10632), .B0(n9886), .B1(n10325), .Y(n8072) );
  NOR2X1TS U7682 ( .A(n10026), .B(n11450), .Y(n7770) );
  NOR2X1TS U7681 ( .A(n11475), .B(n11078), .Y(n7125) );
  OAI22X1TS U7680 ( .A0(n7770), .A1(n12305), .B0(n7125), .B1(n7134), .Y(n8094)
         );
  INVX2TS U8600 ( .A(n7523), .Y(n7890) );
  OAI22X1TS U7679 ( .A0(n7890), .A1(n11486), .B0(n9826), .B1(n7536), .Y(n8095)
         );
  AOI211X1TS U7678 ( .A0(n9885), .A1(n7250), .B0(n8094), .C0(n8095), .Y(n8073)
         );
  NOR2X1TS U8448 ( .A(n10687), .B(n9472), .Y(n7123) );
  AOI22X1TS U7677 ( .A0(n11563), .A1(n8092), .B0(n11533), .B1(n10258), .Y(
        n8086) );
  NOR2X1TS U7676 ( .A(n12114), .B(n11807), .Y(n7898) );
  AOI211X1TS U7674 ( .A0(n10026), .A1(n11534), .B0(n7898), .C0(n8091), .Y(
        n8087) );
  NOR2X1TS U7673 ( .A(n11456), .B(n10018), .Y(n7549) );
  AOI211X1TS U7670 ( .A0(n11480), .A1(n11627), .B0(n8089), .C0(n8090), .Y(
        n8088) );
  AOI211X1TS U7661 ( .A0(n11568), .A1(n11481), .B0(n8082), .C0(n8083), .Y(
        n8079) );
  AOI21X1TS U7658 ( .A0(n12075), .A1(n12463), .B0(n10682), .Y(n8075) );
  INVX2TS U8543 ( .A(n12305), .Y(n8047) );
  AOI22X1TS U7651 ( .A0(n11481), .A1(n10025), .B0(n11443), .B1(n11037), .Y(
        n8066) );
  NOR2X1TS U7650 ( .A(n11159), .B(n11076), .Y(n7766) );
  AOI22X1TS U7648 ( .A0(n11160), .A1(n11082), .B0(n10735), .B1(n7513), .Y(
        n8067) );
  NOR2X1TS U7647 ( .A(n10324), .B(n10058), .Y(n7252) );
  OAI22X1TS U7646 ( .A0(n9806), .A1(n10627), .B0(n7252), .B1(n12095), .Y(n8070) );
  OAI211X1TS U7643 ( .A0(n12561), .A1(n10678), .B0(n7877), .C0(n7870), .Y(
        n8071) );
  AOI211X1TS U7642 ( .A0(n11627), .A1(n10633), .B0(n8070), .C0(n8071), .Y(
        n8068) );
  NOR2X1TS U7639 ( .A(n10329), .B(n11808), .Y(n7894) );
  AOI211X1TS U7637 ( .A0(n11474), .A1(n11563), .B0(n7894), .C0(n8064), .Y(
        n8062) );
  OAI211X1TS U7636 ( .A0(n12561), .A1(n11934), .B0(n8062), .C0(n8063), .Y(
        n8036) );
  OAI22X1TS U7634 ( .A0(n7890), .A1(n10609), .B0(n10681), .B1(n11043), .Y(
        n7360) );
  NOR2X1TS U7632 ( .A(n11160), .B(n11475), .Y(n7880) );
  OAI22X1TS U7628 ( .A0(n12096), .A1(n10678), .B0(n12337), .B1(n12462), .Y(
        n8052) );
  NOR2X1TS U8498 ( .A(n11449), .B(n10258), .Y(n7367) );
  NOR2X1TS U7626 ( .A(n11037), .B(n12089), .Y(n7535) );
  AOI22X1TS U7622 ( .A0(n11443), .A1(n10277), .B0(n9471), .B1(n7753), .Y(n8039) );
  NOR2X1TS U8437 ( .A(n11570), .B(n10058), .Y(n8044) );
  NOR2X1TS U8573 ( .A(n10609), .B(n10005), .Y(n8048) );
  OAI211X1TS U7618 ( .A0(n8044), .A1(n12561), .B0(n8045), .C0(n8046), .Y(n8040) );
  AOI22X1TS U7617 ( .A0(n11444), .A1(n11451), .B0(n11039), .B1(n10320), .Y(
        n8042) );
  OAI211X1TS U7616 ( .A0(n12559), .A1(n10608), .B0(n8042), .C0(n8043), .Y(
        n8041) );
  NOR2X1TS U7615 ( .A(n8040), .B(n8041), .Y(n7506) );
  NOR2X1TS U8227 ( .A(n9602), .B(sa31[7]), .Y(n8468) );
  NOR2X1TS U8080 ( .A(n9865), .B(n11914), .Y(n7835) );
  INVX2TS U8079 ( .A(n7835), .Y(n7487) );
  NOR2X1TS U8224 ( .A(n8467), .B(sa31[3]), .Y(n8463) );
  OAI31X1TS U8077 ( .A0(n11553), .A1(n12362), .A2(n10728), .B0(n12185), .Y(
        n8446) );
  NOR2X1TS U8220 ( .A(n9603), .B(n9373), .Y(n8425) );
  NOR2X1TS U8209 ( .A(n9585), .B(sa31[0]), .Y(n8477) );
  AOI31X1TS U8076 ( .A0(n11521), .A1(n12357), .A2(n10074), .B0(n10029), .Y(
        n8448) );
  NOR2X1TS U8196 ( .A(n9589), .B(sa31[5]), .Y(n8327) );
  AOI211X1TS U8073 ( .A0(n12349), .A1(n11155), .B0(n8448), .C0(n8449), .Y(
        n8447) );
  NOR2X1TS U7610 ( .A(n12143), .B(n11926), .Y(n7667) );
  INVX2TS U8214 ( .A(n8478), .Y(n8443) );
  AOI21X1TS U7609 ( .A0(n11103), .A1(n11920), .B0(n10061), .Y(n7687) );
  NOR2X1TS U7890 ( .A(n10728), .B(n11140), .Y(n7833) );
  NOR2X1TS U7929 ( .A(n11862), .B(n10316), .Y(n7828) );
  OAI211X1TS U7606 ( .A0(n7667), .A1(n11510), .B0(n8033), .C0(n8034), .Y(n8032) );
  AOI211X1TS U7605 ( .A0(n11898), .A1(n12361), .B0(n8031), .C0(n8032), .Y(
        n8015) );
  AOI22X1TS U7604 ( .A0(n7325), .A1(n11616), .B0(n11515), .B1(n10315), .Y(
        n8016) );
  NOR2X1TS U7603 ( .A(n10723), .B(n11107), .Y(n7311) );
  NOR2X1TS U7602 ( .A(n9846), .B(n11921), .Y(n7857) );
  NOR2X1TS U8145 ( .A(n11617), .B(n11138), .Y(n8441) );
  NOR2X1TS U8070 ( .A(n11916), .B(n10315), .Y(n7850) );
  OAI211X1TS U8063 ( .A0(n10711), .A1(n10723), .B0(n8439), .C0(n7684), .Y(
        n8029) );
  NOR2X1TS U7601 ( .A(n9865), .B(n7313), .Y(n7494) );
  AOI22X1TS U8134 ( .A0(n11552), .A1(n12141), .B0(n7315), .B1(n11123), .Y(
        n8464) );
  NOR2X1TS U8128 ( .A(n10661), .B(n10655), .Y(n7821) );
  AOI211X1TS U8126 ( .A0(n12191), .A1(n7686), .B0(n7821), .C0(n8316), .Y(n8465) );
  OAI21X1TS U7596 ( .A0(n12191), .A1(n10729), .B0(n11151), .Y(n8024) );
  NOR2X1TS U7927 ( .A(n10070), .B(n11096), .Y(n7681) );
  NOR2X1TS U7920 ( .A(n10066), .B(n10656), .Y(n8027) );
  AOI211X1TS U7593 ( .A0(n12363), .A1(n11927), .B0(n8027), .C0(n8028), .Y(
        n8026) );
  NOR2X1TS U7891 ( .A(n12357), .B(n10712), .Y(n8013) );
  AOI22X1TS U8190 ( .A0(n11553), .A1(n11515), .B0(n11124), .B1(n7332), .Y(
        n8471) );
  NOR2X1TS U8182 ( .A(n12356), .B(n10648), .Y(n8317) );
  NOR2X1TS U8179 ( .A(n10656), .B(n11610), .Y(n8301) );
  AOI211X1TS U8178 ( .A0(n11144), .A1(n11916), .B0(n8317), .C0(n8301), .Y(
        n8472) );
  OAI21X1TS U8158 ( .A0(n10729), .A1(n11139), .B0(n10282), .Y(n8476) );
  AOI211X1TS U8153 ( .A0(n12634), .A1(n11138), .B0(n8474), .C0(n8475), .Y(
        n8473) );
  OAI211X1TS U7585 ( .A0(n7828), .A1(n11866), .B0(n8011), .C0(n8012), .Y(n7998) );
  OAI22X1TS U7584 ( .A0(n7834), .A1(n11102), .B0(n10030), .B1(n11921), .Y(
        n8005) );
  AOI22X1TS U7582 ( .A0(n12185), .A1(n9543), .B0(n12362), .B1(n12143), .Y(
        n8008) );
  AOI22X1TS U7581 ( .A0(n12183), .A1(n11615), .B0(n12361), .B1(n10281), .Y(
        n8009) );
  AOI211X1TS U7578 ( .A0(n12369), .A1(n7689), .B0(n8005), .C0(n8006), .Y(n7708) );
  AOI22X1TS U7575 ( .A0(n7650), .A1(n7664), .B0(n12617), .B1(n7838), .Y(n8001)
         );
  NOR2X1TS U7574 ( .A(n11527), .B(n10651), .Y(n7816) );
  AOI211X1TS U7572 ( .A0(n10316), .A1(n12632), .B0(n7816), .C0(n8003), .Y(
        n8002) );
  NOR4X1TS U7570 ( .A(n7997), .B(n7477), .C(n7998), .D(n7999), .Y(n1517) );
  INVX2TS U7569 ( .A(n1517), .Y(n1519) );
  AOI31X1TS U8392 ( .A0(n11118), .A1(n11585), .A2(n10094), .B0(n12157), .Y(
        n8541) );
  AOI22X1TS U8380 ( .A0(n11492), .A1(n11504), .B0(n12595), .B1(n8197), .Y(
        n8543) );
  AOI32X1TS U8373 ( .A0(n8543), .A1(n11891), .A2(n10696), .B0(n10356), .B1(
        n8543), .Y(n8542) );
  AOI211X1TS U8372 ( .A0(n9628), .A1(n12470), .B0(n8541), .C0(n8542), .Y(n8536) );
  OAI21X1TS U8365 ( .A0(n10702), .A1(n12135), .B0(n12472), .Y(n8537) );
  OAI32X1TS U8352 ( .A0(n9511), .A1(n8204), .A2(n12596), .B0(n11909), .B1(
        n8204), .Y(n8538) );
  OAI22X1TS U8253 ( .A0(n10093), .A1(n11647), .B0(n11587), .B1(n10050), .Y(
        n8499) );
  OAI32X1TS U8252 ( .A0(n11091), .A1(n8499), .A2(n11945), .B0(n10101), .B1(
        n8499), .Y(n8497) );
  NOR3X1TS U8245 ( .A(n8494), .B(n8390), .C(n8495), .Y(n8492) );
  NOR2X1TS U8244 ( .A(n11193), .B(n10692), .Y(n7275) );
  OAI211X1TS U8241 ( .A0(n7298), .A1(n11951), .B0(n8492), .C0(n8493), .Y(n8227) );
  OAI22X1TS U7863 ( .A0(n11891), .A1(n8270), .B0(n10351), .B1(n12127), .Y(
        n8268) );
  AOI21X1TS U7862 ( .A0(n11646), .A1(n11652), .B0(n11587), .Y(n8269) );
  AOI211X1TS U7861 ( .A0(n10333), .A1(n9531), .B0(n8268), .C0(n8269), .Y(n8267) );
  AOI22X1TS U7857 ( .A0(n11086), .A1(n11093), .B0(n10739), .B1(n7460), .Y(
        n8262) );
  OAI31X1TS U7856 ( .A0(n10702), .A1(n12136), .A2(n9510), .B0(n11580), .Y(
        n8263) );
  OAI211X1TS U7855 ( .A0(n11585), .A1(n11891), .B0(n8262), .C0(n8263), .Y(
        n8241) );
  AOI22X1TS U7852 ( .A0(n11492), .A1(n11910), .B0(n12628), .B1(n12472), .Y(
        n8257) );
  AOI22X1TS U7850 ( .A0(n11194), .A1(n9515), .B0(n12480), .B1(n7593), .Y(n8258) );
  OAI21X1TS U7849 ( .A0(n10638), .A1(n10089), .B0(n10301), .Y(n7612) );
  OAI21X1TS U8259 ( .A0(n10696), .A1(n12127), .B0(n8398), .Y(n8502) );
  AOI21X1TS U8258 ( .A0(n10311), .A1(n12636), .B0(n8502), .Y(n8501) );
  AOI211X1TS U8256 ( .A0(n9629), .A1(n7599), .B0(n8217), .C0(n8500), .Y(n8245)
         );
  OAI22X1TS U7847 ( .A0(n10094), .A1(n10352), .B0(n12157), .B1(n11183), .Y(
        n8251) );
  AOI22X1TS U7845 ( .A0(n12637), .A1(n9628), .B0(n10638), .B1(n10692), .Y(
        n8254) );
  AOI211X1TS U7842 ( .A0(n11499), .A1(n8216), .B0(n8251), .C0(n8252), .Y(n7954) );
  NOR2X1TS U7839 ( .A(n12129), .B(n10749), .Y(n7297) );
  AOI211X1TS U7838 ( .A0(n12179), .A1(n8210), .B0(n8205), .C0(n7297), .Y(n8246) );
  NOR2X1TS U7837 ( .A(n11182), .B(n11645), .Y(n7632) );
  NOR2X1TS U8294 ( .A(n11951), .B(n11165), .Y(n7621) );
  NOR2X1TS U8293 ( .A(n12625), .B(n12478), .Y(n8503) );
  AOI211X1TS U8285 ( .A0(n11172), .A1(n11909), .B0(n7621), .C0(n8517), .Y(
        n8516) );
  OAI211X1TS U8284 ( .A0(n8182), .A1(n10351), .B0(n8363), .C0(n8516), .Y(n8248) );
  AOI22X1TS U7833 ( .A0(n12472), .A1(n11087), .B0(n12179), .B1(n8240), .Y(
        n8229) );
  NOR2X1TS U7832 ( .A(n11170), .B(n12136), .Y(n7585) );
  NOR2X1TS U7987 ( .A(n7629), .B(n11647), .Y(n8239) );
  AOI211X1TS U7829 ( .A0(n11504), .A1(n10311), .B0(n8238), .C0(n8239), .Y(
        n8235) );
  OAI211X1TS U7826 ( .A0(n7459), .A1(n11178), .B0(n8235), .C0(n8236), .Y(n8233) );
  AOI211X1TS U7825 ( .A0(n11194), .A1(n7460), .B0(n8232), .C0(n8233), .Y(n8230) );
  NOR4X1TS U7822 ( .A(n8226), .B(n8227), .C(n7955), .D(n8228), .Y(n1641) );
  INVX2TS U7820 ( .A(n1641), .Y(n1643) );
  INVX2TS U7567 ( .A(n7001), .Y(n6998) );
  AOI22X1TS U8117 ( .A0(n11855), .A1(n12185), .B0(n11139), .B1(n7712), .Y(
        n8457) );
  AOI22X1TS U8115 ( .A0(n12362), .A1(n11516), .B0(n12142), .B1(n10315), .Y(
        n8458) );
  NOR2X1TS U8111 ( .A(n11156), .B(n11097), .Y(n7690) );
  OAI211X1TS U8103 ( .A0(n11866), .A1(n9862), .B0(n7845), .C0(n8321), .Y(n8462) );
  AOI211X1TS U8102 ( .A0(n12190), .A1(n12184), .B0(n8461), .C0(n8462), .Y(
        n8460) );
  NOR2X1TS U8044 ( .A(n11515), .B(n7698), .Y(n7496) );
  OAI22X1TS U7248 ( .A0(n7494), .A1(n11558), .B0(n7496), .B1(n9520), .Y(n7493)
         );
  AOI211X1TS U7247 ( .A0(n11123), .A1(n7491), .B0(n7492), .C0(n7493), .Y(n7470) );
  AOI22X1TS U8062 ( .A0(n11855), .A1(n11926), .B0(n12351), .B1(n11616), .Y(
        n8434) );
  OAI31X1TS U8058 ( .A0(n11861), .A1(n12361), .A2(n10081), .B0(n11958), .Y(
        n8438) );
  AOI211X1TS U8056 ( .A0(n10069), .A1(n12618), .B0(n8436), .C0(n8437), .Y(
        n8435) );
  AOI22X1TS U7363 ( .A0(n11915), .A1(n12184), .B0(n10081), .B1(n11593), .Y(
        n7732) );
  NOR2X1TS U8083 ( .A(n12183), .B(n12143), .Y(n7729) );
  NOR2X1TS U7906 ( .A(n10285), .B(n10713), .Y(n7728) );
  AOI22X1TS U7245 ( .A0(n11896), .A1(n7485), .B0(n12634), .B1(n7487), .Y(n7484) );
  AOI22X1TS U7242 ( .A0(n11898), .A1(n11552), .B0(n10316), .B1(n12617), .Y(
        n7472) );
  AOI22X1TS U8342 ( .A0(n10302), .A1(n12480), .B0(n12178), .B1(n12135), .Y(
        n8532) );
  AOI31X1TS U8339 ( .A0(n11199), .A1(n11585), .A2(n12128), .B0(n11166), .Y(
        n8534) );
  NOR2X1TS U8338 ( .A(n10697), .B(n11199), .Y(n8371) );
  AOI211X1TS U8337 ( .A0(n11580), .A1(n11491), .B0(n8534), .C0(n8371), .Y(
        n8533) );
  AOI211X1TS U8331 ( .A0(n12626), .A1(n11944), .B0(n8415), .C0(n8531), .Y(
        n8530) );
  OAI211X1TS U8327 ( .A0(n10357), .A1(n10749), .B0(n8530), .C0(n8200), .Y(
        n7442) );
  OAI22X1TS U8275 ( .A0(n10347), .A1(n12172), .B0(n8209), .B1(n11177), .Y(
        n8505) );
  OAI211X1TS U8272 ( .A0(n11654), .A1(n10046), .B0(n8510), .C0(n8189), .Y(
        n8508) );
  NOR2X1TS U8316 ( .A(n11498), .B(n10740), .Y(n7963) );
  NOR2X1TS U8271 ( .A(n7986), .B(n11087), .Y(n7587) );
  OAI22X1TS U8270 ( .A0(n7963), .A1(n10086), .B0(n7587), .B1(n10697), .Y(n8509) );
  AOI211X1TS U8269 ( .A0(n12637), .A1(n7610), .B0(n8508), .C0(n8509), .Y(n8507) );
  OAI211X1TS U8267 ( .A0(n12155), .A1(n9877), .B0(n8507), .C0(n8395), .Y(n8506) );
  AOI211X1TS U8266 ( .A0(n10332), .A1(n12596), .B0(n8505), .C0(n8506), .Y(
        n7469) );
  AOI211X1TS U7559 ( .A0(n10691), .A1(n12641), .B0(n7984), .C0(n7985), .Y(
        n7983) );
  OAI211X1TS U7558 ( .A0(n12157), .A1(n11951), .B0(n7982), .C0(n7983), .Y(
        n7981) );
  AOI211X1TS U7557 ( .A0(n8351), .A1(n7979), .B0(n7980), .C0(n7981), .Y(n7977)
         );
  OAI211X1TS U7556 ( .A0(n11176), .A1(n9878), .B0(n7977), .C0(n7978), .Y(n7444) );
  AOI22X1TS U7237 ( .A0(n10301), .A1(n9515), .B0(n11092), .B1(n7460), .Y(n7456) );
  AOI211X1TS U7235 ( .A0(n11491), .A1(n7451), .B0(n7452), .C0(n7453), .Y(n7448) );
  AOI22X1TS U7234 ( .A0(n12637), .A1(n12478), .B0(n12471), .B1(n9510), .Y(
        n7449) );
  OAI211X1TS U7233 ( .A0(n10045), .A1(n10049), .B0(n7448), .C0(n7449), .Y(
        n7445) );
  INVX2TS U7228 ( .A(n7018), .Y(n1282) );
  AOI22X1TS U7555 ( .A0(n10306), .A1(n11579), .B0(n12178), .B1(n12595), .Y(
        n7615) );
  OAI22X1TS U7983 ( .A0(n10046), .A1(n12170), .B0(n11199), .B1(n11641), .Y(
        n8374) );
  NOR2X1TS U7981 ( .A(n8374), .B(n8375), .Y(n7617) );
  AOI22X1TS U7306 ( .A0(n11091), .A1(n9487), .B0(n12473), .B1(n9531), .Y(n7603) );
  AOI211X1TS U7302 ( .A0(n7446), .A1(n7599), .B0(n7600), .C0(n7601), .Y(n7598)
         );
  AOI22X1TS U7988 ( .A0(n11192), .A1(n12136), .B0(n10089), .B1(n12472), .Y(
        n8376) );
  OAI22X1TS U7986 ( .A0(n11118), .A1(n11164), .B0(n11891), .B1(n12129), .Y(
        n8378) );
  AOI211X1TS U7985 ( .A0(n8249), .A1(n9628), .B0(n8239), .C0(n8378), .Y(n8377)
         );
  OAI211X1TS U7984 ( .A0(n8250), .A1(n7989), .B0(n8376), .C0(n8377), .Y(n7265)
         );
  OAI21X1TS U7980 ( .A0(n10745), .A1(n11585), .B0(n8373), .Y(n8372) );
  AOI211X1TS U7979 ( .A0(n10302), .A1(n12627), .B0(n8371), .C0(n8372), .Y(
        n7270) );
  OAI22X1TS U8456 ( .A0(n11932), .A1(n9837), .B0(n12463), .B1(n12306), .Y(
        n7261) );
  NOR2X1TS U8525 ( .A(n11569), .B(n10622), .Y(n7263) );
  AOI211X1TS U7151 ( .A0(n11039), .A1(n7121), .B0(n7261), .C0(n7262), .Y(n7219) );
  NOR2X1TS U8479 ( .A(n10278), .B(n12640), .Y(n7246) );
  AOI22X1TS U7150 ( .A0(n11083), .A1(n10634), .B0(n10026), .B1(n9472), .Y(
        n7255) );
  OAI211X1TS U7149 ( .A0(n12320), .A1(n12101), .B0(n7255), .C0(n7256), .Y(
        n7136) );
  AOI211X1TS U7147 ( .A0(n12313), .A1(n7250), .B0(n7136), .C0(n7251), .Y(n7247) );
  OAI211X1TS U7145 ( .A0(n7246), .A1(n11807), .B0(n7247), .C0(n7248), .Y(n7221) );
  NOR2X1TS U8531 ( .A(n11874), .B(n9817), .Y(n7537) );
  AOI211X1TS U7273 ( .A0(n10058), .A1(n11474), .B0(n7537), .C0(n7538), .Y(
        n7503) );
  NOR2X1TS U7383 ( .A(n10328), .B(n12305), .Y(n7533) );
  OAI22X1TS U7272 ( .A0(n7535), .A1(n10034), .B0(n7263), .B1(n12094), .Y(n7534) );
  AOI211X1TS U7271 ( .A0(n10321), .A1(n12639), .B0(n7533), .C0(n7534), .Y(
        n7530) );
  OAI211X1TS U7270 ( .A0(n11850), .A1(n7569), .B0(n7530), .C0(n7531), .Y(n7098) );
  NOR3X1TS U7471 ( .A(n11039), .B(n11083), .C(n11449), .Y(n7520) );
  OAI22X1TS U7470 ( .A0(n11112), .A1(n11129), .B0(n11849), .B1(n7140), .Y(
        n7529) );
  NOR2X1TS U7476 ( .A(n7880), .B(n11129), .Y(n7524) );
  AOI211X1TS U7267 ( .A0(n10265), .A1(n7523), .B0(n7524), .C0(n7525), .Y(n7522) );
  OAI211X1TS U7266 ( .A0(n7520), .A1(n11806), .B0(n7521), .C0(n7522), .Y(n7504) );
  OAI22X1TS U7265 ( .A0(n12113), .A1(n9838), .B0(n12121), .B1(n12464), .Y(
        n7517) );
  NOR2X1TS U7263 ( .A(n7517), .B(n7518), .Y(n7137) );
  NOR2X1TS U8461 ( .A(n12095), .B(n10628), .Y(n7514) );
  AOI211X1TS U7261 ( .A0(n11565), .A1(n7513), .B0(n7514), .C0(n7515), .Y(n7507) );
  AOI211X1TS U7260 ( .A0(n11535), .A1(n7509), .B0(n7510), .C0(n7511), .Y(n7508) );
  NOR4BX1TS U7258 ( .AN(n7503), .B(n7098), .C(n7504), .D(n7505), .Y(n7223) );
  AOI21X1TS U7143 ( .A0(n10623), .A1(n11481), .B0(n7240), .Y(n7237) );
  OAI211X1TS U7142 ( .A0(n12304), .A1(n12115), .B0(n7236), .C0(n7237), .Y(
        n7232) );
  OAI32X1TS U7141 ( .A0(n7232), .A1(n11473), .A2(n12314), .B0(n11082), .B1(
        n7232), .Y(n7138) );
  AOI22X1TS U7140 ( .A0(n10017), .A1(n12090), .B0(n12639), .B1(n12312), .Y(
        n7224) );
  NOR4BX1TS U7137 ( .AN(n7219), .B(n7220), .C(n7221), .D(n7222), .Y(n6960) );
  OAI22X1TS U8642 ( .A0(n11603), .A1(n10042), .B0(n11771), .B1(n12069), .Y(
        n7189) );
  NOR2X1TS U8711 ( .A(n11879), .B(n11048), .Y(n7191) );
  OAI22X1TS U7121 ( .A0(n7069), .A1(n11770), .B0(n7191), .B1(n11838), .Y(n7190) );
  AOI211X1TS U7120 ( .A0(n11432), .A1(n7067), .B0(n7189), .C0(n7190), .Y(n7147) );
  OAI211X1TS U7118 ( .A0(n11844), .A1(n11794), .B0(n7183), .C0(n7184), .Y(
        n7082) );
  OAI22X1TS U7117 ( .A0(n7180), .A1(n11438), .B0(n9467), .B1(n11421), .Y(n7179) );
  AOI211X1TS U7116 ( .A0(n12553), .A1(n7178), .B0(n7082), .C0(n7179), .Y(n7175) );
  OAI211X1TS U7114 ( .A0(n7174), .A1(n11437), .B0(n7175), .C0(n7176), .Y(n7149) );
  NOR3X1TS U7514 ( .A(n11432), .B(n11463), .C(n11782), .Y(n7432) );
  OAI22X1TS U7513 ( .A0(n11072), .A1(n10298), .B0(n11831), .B1(n10294), .Y(
        n7441) );
  NOR2X1TS U7519 ( .A(n7927), .B(n10297), .Y(n7436) );
  AOI211X1TS U7222 ( .A0(n12455), .A1(n7435), .B0(n7436), .C0(n7437), .Y(n7434) );
  OAI211X1TS U7221 ( .A0(n7432), .A1(n11437), .B0(n7433), .C0(n7434), .Y(n7410) );
  NOR2X1TS U8685 ( .A(n11623), .B(n11050), .Y(n7426) );
  NOR2X1TS U8647 ( .A(n11778), .B(n10618), .Y(n7430) );
  AOI211X1TS U7219 ( .A0(n11885), .A1(n7429), .B0(n7430), .C0(n7431), .Y(n7427) );
  AOI22X1TS U7217 ( .A0(n11790), .A1(n11545), .B0(n11783), .B1(n12550), .Y(
        n7414) );
  NOR2X1TS U8716 ( .A(n11541), .B(n10009), .Y(n7419) );
  NOR2X1TS U7406 ( .A(n10038), .B(n12067), .Y(n7423) );
  OAI211X1TS U7214 ( .A0(n11832), .A1(n11820), .B0(n7420), .C0(n7421), .Y(
        n7044) );
  OAI22X1TS U7212 ( .A0(n11818), .A1(n10042), .B0(n11837), .B1(n11771), .Y(
        n7416) );
  OAI22X1TS U7211 ( .A0(n9810), .A1(n11467), .B0(n11795), .B1(n11539), .Y(
        n7417) );
  NOR2X1TS U7210 ( .A(n7416), .B(n7417), .Y(n7083) );
  AOI21X1TS U7112 ( .A0(n11049), .A1(n11825), .B0(n7168), .Y(n7165) );
  OAI211X1TS U7111 ( .A0(n12070), .A1(n11819), .B0(n7164), .C0(n7165), .Y(
        n7160) );
  NOR4BX1TS U7106 ( .AN(n7147), .B(n7148), .C(n7149), .D(n7150), .Y(n7009) );
  OAI22X1TS U7022 ( .A0(n12656), .A1(n9177), .B0(n7009), .B1(n6960), .Y(n1286)
         );
  NOR2X1TS U8645 ( .A(n11469), .B(n9500), .Y(n7088) );
  OAI21X1TS U7081 ( .A0(n11771), .A1(n11795), .B0(n7091), .Y(n7089) );
  AOI211X1TS U7080 ( .A0(n11783), .A1(n11790), .B0(n7088), .C0(n7089), .Y(
        n7085) );
  OAI22X1TS U7075 ( .A0(n7065), .A1(n9463), .B0(n9797), .B1(n11772), .Y(n7063)
         );
  OAI22X1TS U8671 ( .A0(n9814), .A1(n11764), .B0(n7216), .B1(n9500), .Y(n7064)
         );
  NOR4BX1TS U7074 ( .AN(n7061), .B(n7062), .C(n7063), .D(n7064), .Y(n7048) );
  NOR2X1TS U7412 ( .A(n11818), .B(n9501), .Y(n7053) );
  OAI22X1TS U7206 ( .A0(n7406), .A1(n10037), .B0(n7174), .B1(n12148), .Y(n7398) );
  AOI22X1TS U7204 ( .A0(n12631), .A1(n10614), .B0(n11545), .B1(n12550), .Y(
        n7401) );
  NOR4BX1TS U7202 ( .AN(n7206), .B(n7398), .C(n7399), .D(n7400), .Y(n7058) );
  AOI211X1TS U7071 ( .A0(n7081), .A1(n12629), .B0(n7053), .C0(n7054), .Y(n7049) );
  NOR4X1TS U7069 ( .A(n7043), .B(n7044), .C(n7045), .D(n7046), .Y(n1563) );
  INVX2TS U7068 ( .A(n1563), .Y(n1562) );
  OAI22X1TS U8624 ( .A0(n7786), .A1(n10595), .B0(n8110), .B1(n11830), .Y(n8618) );
  AOI22X1TS U8623 ( .A0(n11824), .A1(n12456), .B0(n9889), .B1(n11633), .Y(
        n8624) );
  AOI32X1TS U8622 ( .A0(n11836), .A1(n8624), .A2(n12327), .B0(n11540), .B1(
        n8624), .Y(n8619) );
  AOI22X1TS U8620 ( .A0(n11884), .A1(n10670), .B0(n11813), .B1(n10590), .Y(
        n8623) );
  AOI32X1TS U8619 ( .A0(n11844), .A1(n8623), .A2(n11427), .B0(n10665), .B1(
        n8623), .Y(n8620) );
  OAI21X1TS U8618 ( .A0(n9890), .A1(n9575), .B0(n12457), .Y(n8622) );
  AOI32X1TS U8617 ( .A0(n12148), .A1(n8622), .A2(n9463), .B0(n11765), .B1(
        n8622), .Y(n8621) );
  OAI22X1TS U7541 ( .A0(n7802), .A1(n11071), .B0(n7798), .B1(n11540), .Y(n7953) );
  AOI31X1TS U7540 ( .A0(n9560), .A1(n7440), .A2(n7797), .B0(n7953), .Y(n7931)
         );
  NOR2X1TS U7538 ( .A(n10269), .B(n10591), .Y(n7787) );
  OAI22X1TS U7537 ( .A0(n7425), .A1(n11439), .B0(n7787), .B1(n10297), .Y(n7951) );
  AOI211X1TS U7536 ( .A0(n11939), .A1(n7395), .B0(n7950), .C0(n7951), .Y(n7932) );
  AOI22X1TS U7535 ( .A0(n11825), .A1(n11621), .B0(n11060), .B1(n12551), .Y(
        n7942) );
  OAI22X1TS U7529 ( .A0(n11819), .A1(n10010), .B0(n10595), .B1(n10664), .Y(
        n7935) );
  AOI22X1TS U7527 ( .A0(n11788), .A1(n11885), .B0(n10013), .B1(n11049), .Y(
        n7939) );
  OAI211X1TS U7526 ( .A0(n7937), .A1(n10297), .B0(n7938), .C0(n7939), .Y(n7936) );
  OAI21X1TS U8681 ( .A0(n11836), .A1(n11842), .B0(n8146), .Y(n8650) );
  AOI22X1TS U8680 ( .A0(n11789), .A1(n11025), .B0(n11634), .B1(n11054), .Y(
        n8652) );
  OAI211X1TS U8678 ( .A0(n10600), .A1(n10009), .B0(n8652), .C0(n8121), .Y(
        n8651) );
  AOI211X1TS U8677 ( .A0(n9890), .A1(n7920), .B0(n8650), .C0(n8651), .Y(n7803)
         );
  OAI211X1TS U7418 ( .A0(n7802), .A1(n7161), .B0(n7803), .C0(n7804), .Y(n7775)
         );
  AOI22X1TS U7414 ( .A0(n11065), .A1(n10289), .B0(n12550), .B1(n7797), .Y(
        n7794) );
  OAI211X1TS U8723 ( .A0(n10665), .A1(n11770), .B0(n7184), .C0(n7091), .Y(
        n8658) );
  OAI32X1TS U8712 ( .A0(n7419), .A1(n11050), .A2(n12455), .B0(n12552), .B1(
        n7419), .Y(n8660) );
  OAI211X1TS U8704 ( .A0(n11837), .A1(n10298), .B0(n8660), .C0(n8661), .Y(
        n8659) );
  AOI211X1TS U8703 ( .A0(n11879), .A1(n11826), .B0(n8658), .C0(n8659), .Y(
        n7777) );
  AOI22X1TS U7407 ( .A0(n11789), .A1(n7788), .B0(n12553), .B1(n7789), .Y(n7778) );
  OAI21X1TS U8211 ( .A0(n11516), .A1(n9870), .B0(n11125), .Y(n8416) );
  OAI22X1TS U8138 ( .A0(n8441), .A1(n10066), .B0(n7321), .B1(n7725), .Y(n8469)
         );
  AOI211X1TS U8137 ( .A0(n12616), .A1(n7836), .B0(n8014), .C0(n8469), .Y(n8417) );
  OAI22X1TS U8099 ( .A0(n11102), .A1(n10062), .B0(n10648), .B1(n10724), .Y(
        n8455) );
  OAI22X1TS U8097 ( .A0(n8004), .A1(n11522), .B0(n10029), .B1(n10337), .Y(
        n8456) );
  NOR2X1TS U8094 ( .A(n9602), .B(n8454), .Y(n7826) );
  AOI22X1TS U8091 ( .A0(n11617), .A1(n7712), .B0(n11928), .B1(n9543), .Y(n8427) );
  NOR2X1TS U8084 ( .A(n8306), .B(n10655), .Y(n7652) );
  OAI22X1TS U8082 ( .A0(n7690), .A1(n11558), .B0(n7729), .B1(n11922), .Y(n8451) );
  AOI211X1TS U8081 ( .A0(n9866), .A1(n8326), .B0(n7652), .C0(n8451), .Y(n8428)
         );
  NOR2X1TS U8052 ( .A(n10343), .B(n10719), .Y(n8322) );
  AOI22X1TS U8051 ( .A0(n12350), .A1(n11097), .B0(n11615), .B1(n10281), .Y(
        n8431) );
  AOI31X1TS U8043 ( .A0(n7496), .A1(n10660), .A2(n10342), .B0(n11511), .Y(
        n8422) );
  AOI211X1TS U8040 ( .A0(n7847), .A1(n7487), .B0(n8422), .C0(n8031), .Y(n8421)
         );
  OAI211X1TS U8038 ( .A0(n7837), .A1(n11599), .B0(n8421), .C0(n8305), .Y(n8420) );
  AOI211X1TS U8037 ( .A0(n11897), .A1(n8340), .B0(n7705), .C0(n8420), .Y(n8419) );
  INVX2TS U8035 ( .A(n9212), .Y(n7028) );
  AOI22X1TS U7066 ( .A0(n6998), .A1(n6927), .B0(n9793), .B1(n7001), .Y(n7041)
         );
  OAI22X1TS U8586 ( .A0(n12114), .A1(n12095), .B0(n10021), .B1(n11485), .Y(
        n8607) );
  OAI22X1TS U8557 ( .A0(n11934), .A1(n12121), .B0(n11848), .B1(n12081), .Y(
        n8609) );
  AOI21X1TS U8552 ( .A0(n11801), .A1(n11044), .B0(n12334), .Y(n8610) );
  OAI211X1TS U8537 ( .A0(n10683), .A1(n12465), .B0(n7256), .C0(n7145), .Y(
        n8592) );
  OAI32X1TS U8527 ( .A0(n7537), .A1(n10622), .A2(n12090), .B0(n7526), .B1(
        n7537), .Y(n8594) );
  OAI22X1TS U8523 ( .A0(n7263), .A1(n10034), .B0(n12096), .B1(n11487), .Y(
        n8596) );
  AOI211X1TS U8519 ( .A0(n11474), .A1(n10622), .B0(n8596), .C0(n8597), .Y(
        n8595) );
  OAI211X1TS U8518 ( .A0(n12119), .A1(n7106), .B0(n8594), .C0(n8595), .Y(n8593) );
  AOI211X1TS U8517 ( .A0(n11569), .A1(n11479), .B0(n8592), .C0(n8593), .Y(
        n7746) );
  OAI22X1TS U8513 ( .A0(n11932), .A1(n11850), .B0(n12096), .B1(n11802), .Y(
        n8587) );
  OAI22X1TS U8511 ( .A0(n9805), .A1(n12115), .B0(n11934), .B1(n10006), .Y(
        n8588) );
  NOR4BX1TS U8504 ( .AN(n8081), .B(n8587), .C(n8588), .D(n8589), .Y(n8586) );
  OAI211X1TS U8501 ( .A0(n10628), .A1(n10022), .B0(n8586), .C0(n7567), .Y(
        n7865) );
  OAI22X1TS U8497 ( .A0(n9825), .A1(n12076), .B0(n7367), .B1(n10053), .Y(n7118) );
  OAI21X1TS U8491 ( .A0(n12122), .A1(n12320), .B0(n8080), .Y(n8583) );
  AOI22X1TS U8490 ( .A0(n11455), .A1(n10604), .B0(n11628), .B1(n10633), .Y(
        n8585) );
  OAI211X1TS U8488 ( .A0(n11044), .A1(n9817), .B0(n8585), .C0(n8055), .Y(n8584) );
  AOI211X1TS U8487 ( .A0(n9885), .A1(n7509), .B0(n8583), .C0(n8584), .Y(n7771)
         );
  AOI211X1TS U8470 ( .A0(n10253), .A1(n11629), .B0(n7510), .C0(n8577), .Y(
        n8566) );
  NOR2X1TS U8467 ( .A(n11443), .B(n11077), .Y(n7365) );
  AOI211X1TS U8463 ( .A0(n11450), .A1(n11473), .B0(n8575), .C0(n8576), .Y(
        n8567) );
  NOR2X1TS U8459 ( .A(n11485), .B(n10053), .Y(n7142) );
  AOI211X1TS U8452 ( .A0(n10320), .A1(n10277), .B0(n8569), .C0(n7887), .Y(
        n8568) );
  AOI22X1TS U8444 ( .A0(n11480), .A1(n7757), .B0(n10057), .B1(n7570), .Y(n8558) );
  NOR2X1TS U8443 ( .A(n11933), .B(n12560), .Y(n8561) );
  AOI211X1TS U8441 ( .A0(n12640), .A1(n11455), .B0(n8561), .C0(n7556), .Y(
        n8559) );
  AOI22X1TS U8440 ( .A0(n11479), .A1(n7124), .B0(n11568), .B1(n10633), .Y(
        n8560) );
  OAI22X1TS U8436 ( .A0(n9830), .A1(n10609), .B0(n8044), .B1(n11848), .Y(n8551) );
  AOI22X1TS U8435 ( .A0(n11479), .A1(n12088), .B0(n9886), .B1(n11627), .Y(
        n8557) );
  AOI22X1TS U8432 ( .A0(n11563), .A1(n10686), .B0(n12639), .B1(n10253), .Y(
        n8556) );
  OAI21X1TS U8430 ( .A0(n9885), .A1(n8047), .B0(n12089), .Y(n8555) );
  AOI32X1TS U8429 ( .A0(n12334), .A1(n8555), .A2(n10006), .B0(n12076), .B1(
        n8555), .Y(n8554) );
  AOI211X1TS U8426 ( .A0(n11450), .A1(n8092), .B0(n8548), .C0(n8549), .Y(n8547) );
  NOR3X1TS U7947 ( .A(n11904), .B(n9589), .C(n9874), .Y(n8334) );
  AOI22X1TS U7943 ( .A0(n12361), .A1(n8326), .B0(n7315), .B1(n8296), .Y(n8337)
         );
  AOI22X1TS U7942 ( .A0(n12369), .A1(n10082), .B0(n12349), .B1(n8340), .Y(
        n8338) );
  AOI211X1TS U7940 ( .A0(n7691), .A1(n7838), .B0(n8334), .C0(n8335), .Y(n7301)
         );
  NOR2X1TS U7939 ( .A(n12355), .B(n11610), .Y(n7740) );
  AOI22X1TS U7934 ( .A0(n12371), .A1(n12190), .B0(n11150), .B1(n7665), .Y(
        n8332) );
  AOI21X1TS U7931 ( .A0(n8327), .A1(n9369), .B0(n12633), .Y(n7317) );
  AOI22X1TS U7930 ( .A0(n10069), .A1(n8326), .B0(n11146), .B1(n9542), .Y(n8324) );
  AOI22X1TS U7925 ( .A0(n12141), .A1(n7485), .B0(n11928), .B1(n7330), .Y(n8325) );
  AOI211X1TS U7923 ( .A0(n7325), .A1(n7836), .B0(n7652), .C0(n8323), .Y(n8307)
         );
  AOI211X1TS U7919 ( .A0(n11616), .A1(n11517), .B0(n8027), .C0(n8322), .Y(
        n8314) );
  OAI211X1TS U7914 ( .A0(n7333), .A1(n10652), .B0(n8314), .C0(n8315), .Y(n7679) );
  OAI22X1TS U7913 ( .A0(n10286), .A1(n10343), .B0(n11599), .B1(n10652), .Y(
        n8309) );
  AOI211X1TS U7903 ( .A0(n12489), .A1(n12190), .B0(n7728), .C0(n8303), .Y(
        n7683) );
  OAI32X1TS U7894 ( .A0(n8295), .A1(n12350), .A2(n11926), .B0(n7716), .B1(
        n8295), .Y(n8294) );
  OAI211X1TS U7892 ( .A0(n10706), .A1(n7733), .B0(n8294), .C0(n7482), .Y(n7646) );
  OAI211X1TS U7887 ( .A0(n7833), .A1(n11610), .B0(n8292), .C0(n8293), .Y(n8291) );
  AOI211X1TS U7886 ( .A0(n11144), .A1(n12189), .B0(n8013), .C0(n8291), .Y(
        n7307) );
  OAI211X1TS U7878 ( .A0(n11609), .A1(n11597), .B0(n8284), .C0(n8285), .Y(
        n8283) );
  AOI21X1TS U7877 ( .A0(n11897), .A1(n11615), .B0(n8283), .Y(n7319) );
  OAI211X1TS U7872 ( .A0(n12355), .A1(n10030), .B0(n8279), .C0(n8280), .Y(
        n7653) );
  INVX2TS U7867 ( .A(n1515), .Y(n1516) );
  OAI22X1TS U7061 ( .A0(n7037), .A1(n12736), .B0(n12682), .B1(n7038), .Y(N116)
         );
  NOR2X1TS U7280 ( .A(n10006), .B(n12462), .Y(n7353) );
  AOI22X1TS U7277 ( .A0(n10258), .A1(n11077), .B0(n10325), .B1(n12314), .Y(
        n7543) );
  OAI22X1TS U7201 ( .A0(n9798), .A1(n10294), .B0(n7174), .B1(n12327), .Y(n7373) );
  NOR2X1TS U8650 ( .A(n10036), .B(n9617), .Y(n7215) );
  AOI21X1TS U7195 ( .A0(n11061), .A1(n10591), .B0(n7383), .Y(n7382) );
  INVX2TS U7190 ( .A(n9181), .Y(n7019) );
  INVX2TS U7256 ( .A(n9160), .Y(n6972) );
  OAI22X1TS U7038 ( .A0(n9160), .A1(n9182), .B0(n7019), .B1(n6972), .Y(n1304)
         );
  INVX2TS U7037 ( .A(n1304), .Y(n1303) );
  OAI22X1TS U7134 ( .A0(n7216), .A1(n11439), .B0(n11072), .B1(n7158), .Y(n7212) );
  AOI22X1TS U7523 ( .A0(n11884), .A1(n10269), .B0(n10590), .B1(n11546), .Y(
        n7921) );
  AOI211X1TS U7516 ( .A0(n11033), .A1(n7925), .B0(n7436), .C0(n7926), .Y(n7923) );
  OAI22X1TS U7131 ( .A0(n7065), .A1(n9810), .B0(n9813), .B1(n11427), .Y(n7201)
         );
  OAI22X1TS U8697 ( .A0(n9797), .A1(n11820), .B0(n11605), .B1(n9463), .Y(n8655) );
  NOR4BX1TS U8690 ( .AN(n8147), .B(n8654), .C(n8655), .D(n8656), .Y(n8653) );
  OAI211X1TS U8687 ( .A0(n10617), .A1(n7940), .B0(n8653), .C0(n7389), .Y(n7911) );
  AOI21X1TS U8670 ( .A0(n11634), .A1(n10590), .B0(n7064), .Y(n8647) );
  OAI31X1TS U8656 ( .A0(n11826), .A1(n9575), .A2(n7214), .B0(n12631), .Y(n8643) );
  AOI22X1TS U8651 ( .A0(n11059), .A1(n11055), .B0(n10013), .B1(n12457), .Y(
        n8632) );
  AOI211X1TS U8638 ( .A0(n10673), .A1(n10274), .B0(n8635), .C0(n7934), .Y(
        n8634) );
  OAI22X1TS U7498 ( .A0(n7770), .A1(n11114), .B0(n7766), .B1(n11872), .Y(n7906) );
  AOI31X1TS U7497 ( .A0(n9555), .A1(n7528), .A2(n7765), .B0(n7906), .Y(n7884)
         );
  NOR2X1TS U7495 ( .A(n10017), .B(n10254), .Y(n7755) );
  OAI22X1TS U7494 ( .A0(n7535), .A1(n11807), .B0(n7755), .B1(n11129), .Y(n7904) );
  AOI211X1TS U7493 ( .A0(n11159), .A1(n7564), .B0(n7903), .C0(n7904), .Y(n7885) );
  AOI22X1TS U7492 ( .A0(n11480), .A1(n10734), .B0(n10025), .B1(n12313), .Y(
        n7895) );
  OAI22X1TS U7486 ( .A0(n12113), .A1(n9818), .B0(n10608), .B1(n10682), .Y(
        n7888) );
  AOI22X1TS U7485 ( .A0(n11565), .A1(n7253), .B0(n12638), .B1(n11475), .Y(
        n7891) );
  AOI22X1TS U7484 ( .A0(n11456), .A1(n11564), .B0(n9471), .B1(n10623), .Y(
        n7892) );
  OAI211X1TS U7483 ( .A0(n7890), .A1(n11128), .B0(n7891), .C0(n7892), .Y(n7889) );
  AOI21X1TS U7393 ( .A0(n11850), .A1(n11806), .B0(n12076), .Y(n7759) );
  OAI22X1TS U7392 ( .A0(n12115), .A1(n12561), .B0(n11872), .B1(n12336), .Y(
        n7760) );
  AOI22X1TS U7391 ( .A0(n11534), .A1(n10057), .B0(n12312), .B1(n7765), .Y(
        n7762) );
  NOR2X1TS U7389 ( .A(n12113), .B(n10054), .Y(n7107) );
  AOI211X1TS U7388 ( .A0(n10325), .A1(n10687), .B0(n7764), .C0(n7107), .Y(
        n7763) );
  OAI211X1TS U7387 ( .A0(n9838), .A1(n12320), .B0(n7762), .C0(n7763), .Y(n7761) );
  OAI22X1TS U7029 ( .A0(n7013), .A1(n12737), .B0(n12683), .B1(n7014), .Y(N129)
         );
  NOR2X1TS U4760 ( .A(n11290), .B(n11400), .Y(n4134) );
  NOR2X1TS U4693 ( .A(n11236), .B(n11314), .Y(n4135) );
  NOR2X1TS U4773 ( .A(n4439), .B(n5038), .Y(n4466) );
  NOR2X1TS U3840 ( .A(n9150), .B(n12427), .Y(n4136) );
  NOR4BX1TS U3617 ( .AN(n4133), .B(n4134), .C(n4135), .D(n4136), .Y(n4124) );
  NOR2X1TS U4829 ( .A(sa22[0]), .B(n9446), .Y(n5043) );
  OAI22X1TS U3616 ( .A0(n9147), .A1(n12397), .B0(n9150), .B1(n10383), .Y(n4129) );
  INVX2TS U4816 ( .A(n9248), .Y(n4117) );
  OAI32X1TS U3615 ( .A0(n4129), .A1(n11278), .A2(n11393), .B0(n11725), .B1(
        n4129), .Y(n4125) );
  NOR2X1TS U3614 ( .A(n10464), .B(n12395), .Y(n3881) );
  NOR2X1TS U4801 ( .A(n12501), .B(n10828), .Y(n4128) );
  OAI22X1TS U3613 ( .A0(n4128), .A1(n10388), .B0(n10893), .B1(n11238), .Y(
        n4127) );
  AOI211X1TS U3612 ( .A0(n9642), .A1(n12229), .B0(n3881), .C0(n4127), .Y(n4126) );
  AOI22X1TS U4060 ( .A0(n10887), .A1(n4454), .B0(n10442), .B1(n11731), .Y(
        n4687) );
  NOR2X1TS U4761 ( .A(n9147), .B(n10471), .Y(n4689) );
  NOR2X1TS U4723 ( .A(n10131), .B(n10467), .Y(n4690) );
  OAI211X1TS U4058 ( .A0(n10117), .A1(n10464), .B0(n4687), .C0(n4688), .Y(
        n4686) );
  OAI211X1TS U4055 ( .A0(n10822), .A1(n10472), .B0(n4684), .C0(n4191), .Y(
        n3778) );
  NOR2X1TS U4087 ( .A(n10381), .B(n11315), .Y(n4708) );
  NOR2X1TS U4086 ( .A(n9147), .B(n11236), .Y(n4453) );
  OAI211X1TS U4078 ( .A0(n4705), .A1(n10468), .B0(n4706), .C0(n4707), .Y(n3779) );
  NOR2X1TS U4758 ( .A(n9911), .B(n12395), .Y(n3798) );
  NOR2X1TS U4041 ( .A(n10127), .B(n11732), .Y(n3768) );
  AOI22X1TS U3437 ( .A0(n11286), .A1(n3791), .B0(n12215), .B1(n3796), .Y(n3782) );
  AOI22X1TS U3436 ( .A0(n11727), .A1(n3791), .B0(n9909), .B1(n9114), .Y(n3783)
         );
  NOR2X1TS U4727 ( .A(n11308), .B(n11985), .Y(n4202) );
  NOR2X1TS U4703 ( .A(n4202), .B(n4221), .Y(n3786) );
  NOR2X1TS U4738 ( .A(n12578), .B(n12214), .Y(n3788) );
  NOR2X1TS U3866 ( .A(n10476), .B(n4466), .Y(n3589) );
  AOI211X1TS U3434 ( .A0(n12246), .A1(n3785), .B0(n3786), .C0(n3787), .Y(n3784) );
  NOR2X1TS U4737 ( .A(n12216), .B(n10443), .Y(n4204) );
  NOR2X1TS U4710 ( .A(n10408), .B(n11322), .Y(n4704) );
  OAI32X1TS U4073 ( .A0(n4699), .A1(n11726), .A2(n3590), .B0(n10887), .B1(
        n4699), .Y(n3740) );
  OAI211X1TS U4096 ( .A0(n11399), .A1(n11296), .B0(n4721), .C0(n4722), .Y(
        n4714) );
  NOR2X1TS U4095 ( .A(n9911), .B(n12430), .Y(n4452) );
  OAI211X1TS U4092 ( .A0(n12397), .A1(n10132), .B0(n4719), .C0(n3886), .Y(
        n4715) );
  AOI22X1TS U4090 ( .A0(n12244), .A1(n11732), .B0(n10780), .B1(n3796), .Y(
        n4717) );
  OAI21X1TS U4718 ( .A0(n12053), .A1(n12215), .B0(n9909), .Y(n4718) );
  OAI211X1TS U4089 ( .A0(n11315), .A1(n11995), .B0(n4717), .C0(n4718), .Y(
        n4716) );
  NOR3X1TS U4088 ( .A(n4714), .B(n4715), .C(n4716), .Y(n3741) );
  NOR2X1TS U4696 ( .A(n11727), .B(n10778), .Y(n3773) );
  NOR2X1TS U3430 ( .A(n10127), .B(n11309), .Y(n3591) );
  NOR2X1TS U4724 ( .A(n10437), .B(n11297), .Y(n3765) );
  NOR2X1TS U4702 ( .A(n9662), .B(n9672), .Y(n4110) );
  NOR4BX1TS U3603 ( .AN(n4109), .B(n4110), .C(n4111), .D(n4112), .Y(n3747) );
  NOR2X1TS U3678 ( .A(n10823), .B(n11237), .Y(n3754) );
  INVX2TS U3418 ( .A(n9163), .Y(n3394) );
  NOR2X1TS U4565 ( .A(n11338), .B(n11412), .Y(n4078) );
  NOR2X1TS U4498 ( .A(n11242), .B(n11363), .Y(n4079) );
  NOR2X1TS U4578 ( .A(n4399), .B(n4980), .Y(n4426) );
  NOR2X1TS U3804 ( .A(n9138), .B(n12444), .Y(n4080) );
  NOR4BX1TS U3584 ( .AN(n4077), .B(n4078), .C(n4079), .D(n4080), .Y(n4068) );
  NOR2X1TS U4634 ( .A(n9828), .B(n9132), .Y(n4985) );
  OAI22X1TS U3583 ( .A0(n9135), .A1(n12403), .B0(n9138), .B1(n10392), .Y(n4073) );
  INVX2TS U4621 ( .A(n9240), .Y(n4061) );
  OAI32X1TS U3582 ( .A0(n4073), .A1(n11328), .A2(n11405), .B0(n11745), .B1(
        n4073), .Y(n4069) );
  NOR2X1TS U3581 ( .A(n10482), .B(n12406), .Y(n3856) );
  NOR2X1TS U4606 ( .A(n12516), .B(n10854), .Y(n4072) );
  OAI22X1TS U3580 ( .A0(n4072), .A1(n10399), .B0(n10910), .B1(n11243), .Y(
        n4071) );
  INVX2TS U4509 ( .A(n12522), .Y(n4177) );
  AOI22X1TS U3985 ( .A0(n10905), .A1(n4414), .B0(n10451), .B1(n11749), .Y(
        n4615) );
  NOR2X1TS U4566 ( .A(n9135), .B(n10489), .Y(n4617) );
  NOR2X1TS U4528 ( .A(n10139), .B(n10485), .Y(n4618) );
  OAI211X1TS U3983 ( .A0(n10110), .A1(n10481), .B0(n4615), .C0(n4616), .Y(
        n4614) );
  OAI211X1TS U3980 ( .A0(n10848), .A1(n10489), .B0(n4612), .C0(n4147), .Y(
        n3712) );
  NOR2X1TS U4011 ( .A(n9135), .B(n11242), .Y(n4413) );
  NOR2X1TS U4563 ( .A(n9915), .B(n12403), .Y(n3732) );
  NOR2X1TS U3966 ( .A(n10135), .B(n11750), .Y(n3702) );
  AOI22X1TS U3412 ( .A0(n11333), .A1(n3725), .B0(n12221), .B1(n3730), .Y(n3716) );
  AOI22X1TS U3411 ( .A0(n11743), .A1(n3725), .B0(n9905), .B1(n9106), .Y(n3717)
         );
  NOR2X1TS U4532 ( .A(n11356), .B(n12000), .Y(n4158) );
  NOR2X1TS U4508 ( .A(n4158), .B(n4177), .Y(n3720) );
  NOR2X1TS U4543 ( .A(n12585), .B(n12222), .Y(n3722) );
  NOR2X1TS U3830 ( .A(n10494), .B(n4426), .Y(n3550) );
  AOI211X1TS U3409 ( .A0(n12270), .A1(n3719), .B0(n3720), .C0(n3721), .Y(n3718) );
  NOR2X1TS U4542 ( .A(n12223), .B(n10450), .Y(n4160) );
  NOR2X1TS U4515 ( .A(n10404), .B(n11368), .Y(n4632) );
  OAI32X1TS U3998 ( .A0(n4627), .A1(n11744), .A2(n12060), .B0(n10905), .B1(
        n4627), .Y(n3674) );
  OAI211X1TS U4021 ( .A0(n11411), .A1(n11345), .B0(n4649), .C0(n4650), .Y(
        n4642) );
  NOR2X1TS U4020 ( .A(n9915), .B(n12445), .Y(n4412) );
  OAI211X1TS U4017 ( .A0(n12405), .A1(n10140), .B0(n4647), .C0(n3861), .Y(
        n4643) );
  AOI22X1TS U4015 ( .A0(n12267), .A1(n11750), .B0(n10766), .B1(n3730), .Y(
        n4645) );
  OAI21X1TS U4523 ( .A0(n12060), .A1(n3701), .B0(n9906), .Y(n4646) );
  OAI211X1TS U4014 ( .A0(n11363), .A1(n12010), .B0(n4645), .C0(n4646), .Y(
        n4644) );
  NOR3X1TS U4013 ( .A(n4642), .B(n4643), .C(n4644), .Y(n3675) );
  NOR2X1TS U4501 ( .A(n11743), .B(n10767), .Y(n3707) );
  NOR2X1TS U3405 ( .A(n10135), .B(n11357), .Y(n3552) );
  NOR2X1TS U4529 ( .A(n10446), .B(n11345), .Y(n3699) );
  NOR2X1TS U4507 ( .A(n9666), .B(n9668), .Y(n4054) );
  OAI22X1TS U3575 ( .A0(n11261), .A1(n10849), .B0(n10424), .B1(n10105), .Y(
        n4055) );
  NOR4BX1TS U3570 ( .AN(n4053), .B(n4054), .C(n4055), .D(n4056), .Y(n3681) );
  NOR2X1TS U3650 ( .A(n10848), .B(n11242), .Y(n3688) );
  NOR2X1TS U5044 ( .A(n10313), .B(n4515), .Y(n5103) );
  NOR2X1TS U5015 ( .A(n11163), .B(n9208), .Y(n4517) );
  AOI22X1TS U4276 ( .A0(n10391), .A1(n12620), .B0(n10812), .B1(n11248), .Y(
        n4842) );
  NOR2X1TS U5034 ( .A(n10319), .B(sa00[5]), .Y(n5092) );
  INVX2TS U5048 ( .A(n5111), .Y(n4475) );
  INVX2TS U4927 ( .A(n9640), .Y(n4841) );
  INVX2TS U4958 ( .A(n9200), .Y(n4334) );
  INVX2TS U5038 ( .A(n9682), .Y(n4840) );
  NOR2X1TS U4271 ( .A(n10803), .B(n10411), .Y(n4503) );
  NOR2X1TS U4934 ( .A(n11702), .B(n12621), .Y(n3953) );
  AOI211X1TS U4266 ( .A0(n11376), .A1(n9680), .B0(n4553), .C0(n4868), .Y(n4844) );
  NOR2X1TS U4264 ( .A(n9901), .B(n12022), .Y(n4497) );
  INVX2TS U5021 ( .A(n9196), .Y(n3947) );
  NOR2X1TS U4261 ( .A(n10860), .B(n10865), .Y(n4486) );
  AOI211X1TS U4260 ( .A0(n10134), .A1(n10415), .B0(n4866), .C0(n4486), .Y(
        n4864) );
  OAI211X1TS U4259 ( .A0(n12567), .A1(n10859), .B0(n4864), .C0(n4865), .Y(
        n4863) );
  OAI32X1TS U4258 ( .A0(n4863), .A1(n12200), .A2(n9687), .B0(n11214), .B1(
        n4863), .Y(n4862) );
  OAI211X1TS U4257 ( .A0(n12572), .A1(n9673), .B0(n4861), .C0(n4862), .Y(n4524) );
  NOR2X1TS U4923 ( .A(n12200), .B(n10148), .Y(n4856) );
  NOR2X1TS U4246 ( .A(n10137), .B(n12031), .Y(n3639) );
  NOR2X1TS U4938 ( .A(n12619), .B(n11250), .Y(n4833) );
  INVX2TS U4937 ( .A(n4833), .Y(n4502) );
  AOI22X1TS U4244 ( .A0(n9690), .A1(n4502), .B0(n10116), .B1(n4306), .Y(n4851)
         );
  NOR2X1TS U4237 ( .A(n10797), .B(n11212), .Y(n4509) );
  NOR2X1TS U4235 ( .A(n9690), .B(n4841), .Y(n3647) );
  NOR2X1TS U4869 ( .A(n10798), .B(n10803), .Y(n4834) );
  OAI22X1TS U4229 ( .A0(n4833), .A1(n12382), .B0(n4834), .B1(n10861), .Y(n4826) );
  OAI22X1TS U4228 ( .A0(n12492), .A1(n12411), .B0(n3954), .B1(n9670), .Y(n4827) );
  AOI21X1TS U4227 ( .A0(n12567), .A1(n11755), .B0(n10775), .Y(n4828) );
  NOR2X1TS U4901 ( .A(n10143), .B(n11380), .Y(n4832) );
  NOR2X1TS U4225 ( .A(n10865), .B(n11714), .Y(n4498) );
  OAI211X1TS U4223 ( .A0(n12538), .A1(n12207), .B0(n4830), .C0(n4831), .Y(
        n4829) );
  NOR2X1TS U4953 ( .A(n10872), .B(n9674), .Y(n4824) );
  INVX2TS U4220 ( .A(n4300), .Y(n3914) );
  NOR2X1TS U4464 ( .A(n4282), .B(n10748), .Y(n4742) );
  NOR2X1TS U4462 ( .A(n9229), .B(n10368), .Y(n4938) );
  NOR2X1TS U4455 ( .A(n9895), .B(n10752), .Y(n4921) );
  AOI22X1TS U4452 ( .A0(n10926), .A1(n10122), .B0(n11219), .B1(n11274), .Y(
        n4904) );
  NOR2X1TS U4433 ( .A(n10120), .B(n9664), .Y(n4732) );
  INVX2TS U4422 ( .A(n9657), .Y(n4903) );
  AOI22X1TS U4416 ( .A0(n11266), .A1(n4900), .B0(n12072), .B1(n11274), .Y(
        n4936) );
  NOR2X1TS U4409 ( .A(n10945), .B(n12277), .Y(n4754) );
  NOR2X1TS U4406 ( .A(n10163), .B(n10402), .Y(n4772) );
  OAI22X1TS U4396 ( .A0(n3837), .A1(n12549), .B0(n12390), .B1(n10123), .Y(
        n4932) );
  AOI211X1TS U4395 ( .A0(n10386), .A1(n11810), .B0(n4364), .C0(n4932), .Y(
        n4906) );
  AOI22X1TS U4393 ( .A0(n10881), .A1(n11792), .B0(n11218), .B1(n11266), .Y(
        n4926) );
  NOR2X1TS U4385 ( .A(n10754), .B(n10922), .Y(n4263) );
  INVX2TS U4383 ( .A(n9225), .Y(n3830) );
  OAI32X1TS U4372 ( .A0(n4924), .A1(n9180), .A2(n12376), .B0(n11798), .B1(
        n4924), .Y(n4923) );
  OAI211X1TS U4369 ( .A0(n12389), .A1(n10755), .B0(n4923), .C0(n4760), .Y(
        n4339) );
  NOR2X1TS U4366 ( .A(n9917), .B(n10126), .Y(n3615) );
  INVX2TS U4365 ( .A(n3615), .Y(n4358) );
  AOI22X1TS U4364 ( .A0(n11797), .A1(n10800), .B0(n11273), .B1(n4358), .Y(
        n4912) );
  NOR2X1TS U4362 ( .A(n12282), .B(n10921), .Y(n4731) );
  OAI32X1TS U4360 ( .A0(n4731), .A1(n9903), .A2(n12074), .B0(n10786), .B1(
        n4731), .Y(n4913) );
  OAI21X1TS U4355 ( .A0(n10927), .A1(n10430), .B0(n11219), .Y(n4919) );
  AOI32X1TS U4354 ( .A0(n10758), .A1(n4919), .A2(n9660), .B0(n12284), .B1(
        n4919), .Y(n4917) );
  AOI211X1TS U4351 ( .A0(n10434), .A1(n4916), .B0(n4917), .C0(n4918), .Y(n4914) );
  NOR2X1TS U4347 ( .A(n11220), .B(n10122), .Y(n4261) );
  AOI22X1TS U4342 ( .A0(n10785), .A1(n4784), .B0(n10125), .B1(n4022), .Y(n4911) );
  NOR2X1TS U4328 ( .A(n10786), .B(n10883), .Y(n3517) );
  OAI211X1TS U4323 ( .A0(n4276), .A1(n10763), .B0(n4898), .C0(n4899), .Y(n4877) );
  NOR2X1TS U4320 ( .A(n11787), .B(n9933), .Y(n4744) );
  OAI22X1TS U4319 ( .A0(n4261), .A1(n9908), .B0(n4744), .B1(n10754), .Y(n4892)
         );
  OAI22X1TS U4318 ( .A0(n11709), .A1(n12037), .B0(n10795), .B1(n10939), .Y(
        n4893) );
  AOI21X1TS U4317 ( .A0(n12390), .A1(n11805), .B0(n10119), .Y(n4894) );
  NOR2X1TS U4316 ( .A(n10152), .B(n10944), .Y(n4770) );
  NOR2X1TS U4315 ( .A(n10922), .B(n10763), .Y(n4252) );
  OAI211X1TS U4312 ( .A0(n10757), .A1(n12066), .B0(n4896), .C0(n4897), .Y(
        n4895) );
  NOR2X1TS U4309 ( .A(n10499), .B(n9661), .Y(n4778) );
  NOR2X1TS U4308 ( .A(n11219), .B(n11785), .Y(n3616) );
  NOR2X1TS U4304 ( .A(n10944), .B(n4243), .Y(n4791) );
  NOR2X1TS U4302 ( .A(n10498), .B(n10164), .Y(n4775) );
  NOR2X1TS U4301 ( .A(n10756), .B(n10503), .Y(n4787) );
  AOI211X1TS U4300 ( .A0(n10433), .A1(n4781), .B0(n4775), .C0(n4787), .Y(n4889) );
  OAI211X1TS U4298 ( .A0(n9929), .A1(n9907), .B0(n4889), .C0(n4262), .Y(n4888)
         );
  AOI211X1TS U4297 ( .A0(n10160), .A1(n10129), .B0(n4791), .C0(n4888), .Y(
        n4359) );
  NOR2X1TS U4296 ( .A(n12378), .B(n10932), .Y(n4247) );
  OAI21X1TS U4289 ( .A0(n11417), .A1(n9918), .B0(n11268), .Y(n4887) );
  OAI211X1TS U4287 ( .A0(n11804), .A1(n12284), .B0(n4887), .C0(n3997), .Y(
        n4884) );
  OAI21X1TS U4286 ( .A0(n10369), .A1(n11786), .B0(n10934), .Y(n4886) );
  OAI211X1TS U4284 ( .A0(n12038), .A1(n10788), .B0(n4886), .C0(n3624), .Y(
        n4885) );
  OAI21X1TS U4282 ( .A0(n10375), .A1(n10784), .B0(n11811), .Y(n4880) );
  AOI22X1TS U4280 ( .A0(n11417), .A1(n3620), .B0(n10429), .B1(n9917), .Y(n4881) );
  OAI22X1TS U3363 ( .A0(n3589), .A1(n10463), .B0(n3591), .B1(n9911), .Y(n3588)
         );
  OAI211X1TS U3361 ( .A0(n3582), .A1(n12429), .B0(n3584), .C0(n3585), .Y(n3559) );
  AOI22X1TS U3360 ( .A0(n12246), .A1(n10888), .B0(n12236), .B1(n3581), .Y(
        n3576) );
  OAI211X1TS U3359 ( .A0(n10895), .A1(n10468), .B0(n3576), .C0(n3577), .Y(
        n3560) );
  OAI22X1TS U4042 ( .A0(n3788), .A1(n11254), .B0(n4667), .B1(n10383), .Y(n4661) );
  OAI22X1TS U4040 ( .A0(n3768), .A1(n11303), .B0(n9161), .B1(n12396), .Y(n4662) );
  AOI22X1TS U4037 ( .A0(n11726), .A1(n9643), .B0(n10828), .B1(n12507), .Y(
        n4665) );
  AOI32X1TS U4036 ( .A0(n4665), .A1(n11398), .A2(n11304), .B0(n10118), .B1(
        n4665), .Y(n4664) );
  NOR2X1TS U4052 ( .A(n10420), .B(n10471), .Y(n4446) );
  NOR2X1TS U4839 ( .A(n3803), .B(n10372), .Y(n4678) );
  OAI21X1TS U4051 ( .A0(n11725), .A1(n11224), .B0(n12236), .Y(n4679) );
  AOI22X1TS U4050 ( .A0(n10804), .A1(n10828), .B0(n11727), .B1(n10774), .Y(
        n4680) );
  AOI211X1TS U4048 ( .A0(n11320), .A1(n10889), .B0(n4446), .C0(n4677), .Y(
        n3563) );
  NOR2X1TS U4757 ( .A(n10118), .B(n11316), .Y(n4089) );
  OAI22X1TS U3597 ( .A0(n4099), .A1(n9912), .B0(n11302), .B1(n11237), .Y(n4090) );
  AOI21X1TS U3594 ( .A0(n11302), .A1(n10463), .B0(n10816), .Y(n4096) );
  OAI32X1TS U3593 ( .A0(n4096), .A1(n11309), .A2(n12237), .B0(n10804), .B1(
        n4096), .Y(n4093) );
  INVX2TS U3323 ( .A(n9092), .Y(n1596) );
  NOR2X1TS U6643 ( .A(n11311), .B(n11217), .Y(n5934) );
  NOR2X1TS U6576 ( .A(n11389), .B(n11287), .Y(n5935) );
  NOR2X1TS U6656 ( .A(n6242), .B(n6837), .Y(n6269) );
  NOR2X1TS U5722 ( .A(n9349), .B(n12399), .Y(n5936) );
  NOR4BX1TS U5500 ( .AN(n5933), .B(n5934), .C(n5935), .D(n5936), .Y(n5924) );
  NOR2X1TS U6712 ( .A(n9880), .B(n9343), .Y(n6842) );
  OAI22X1TS U5499 ( .A0(n9346), .A1(n12423), .B0(n9349), .B1(n10542), .Y(n5929) );
  INVX2TS U6699 ( .A(n9444), .Y(n5917) );
  OAI32X1TS U5498 ( .A0(n5929), .A1(n11325), .A2(n11222), .B0(n11705), .B1(
        n5929), .Y(n5925) );
  NOR2X1TS U5497 ( .A(n10453), .B(n12426), .Y(n5711) );
  NOR2X1TS U6684 ( .A(n12527), .B(n10912), .Y(n5928) );
  OAI22X1TS U5496 ( .A0(n5928), .A1(n10536), .B0(n10873), .B1(n11390), .Y(
        n5927) );
  INVX2TS U6587 ( .A(n12518), .Y(n6131) );
  AOI22X1TS U5943 ( .A0(n10878), .A1(n6257), .B0(n10465), .B1(n11698), .Y(
        n6487) );
  NOR2X1TS U6644 ( .A(n9346), .B(n10444), .Y(n6489) );
  NOR2X1TS U6606 ( .A(n10165), .B(n10448), .Y(n6490) );
  OAI211X1TS U5941 ( .A0(n10221), .A1(n10453), .B0(n6487), .C0(n6488), .Y(
        n6486) );
  OAI211X1TS U5938 ( .A0(n10919), .A1(n10444), .B0(n6484), .C0(n6101), .Y(
        n5533) );
  NOR2X1TS U5969 ( .A(n9346), .B(n11389), .Y(n6256) );
  NOR2X1TS U6641 ( .A(n9949), .B(n12423), .Y(n5553) );
  NOR2X1TS U5924 ( .A(n10169), .B(n11699), .Y(n5523) );
  AOI22X1TS U5308 ( .A0(n11318), .A1(n5546), .B0(n12271), .B1(n5551), .Y(n5537) );
  AOI22X1TS U5307 ( .A0(n11706), .A1(n5546), .B0(n9961), .B1(n9307), .Y(n5538)
         );
  NOR2X1TS U6610 ( .A(n11293), .B(n12047), .Y(n6112) );
  NOR2X1TS U6586 ( .A(n6112), .B(n6131), .Y(n5541) );
  NOR2X1TS U6621 ( .A(n12589), .B(n12272), .Y(n5543) );
  NOR2X1TS U5748 ( .A(n10440), .B(n6269), .Y(n5387) );
  AOI211X1TS U5305 ( .A0(n12242), .A1(n5540), .B0(n5541), .C0(n5542), .Y(n5539) );
  NOR2X1TS U6620 ( .A(n12273), .B(n10466), .Y(n6114) );
  NOR2X1TS U6593 ( .A(n10585), .B(n11281), .Y(n6504) );
  OAI32X1TS U5956 ( .A0(n6499), .A1(n11705), .A2(n11972), .B0(n10880), .B1(
        n6499), .Y(n5495) );
  OAI211X1TS U5979 ( .A0(n11216), .A1(n11306), .B0(n6521), .C0(n6522), .Y(
        n6514) );
  NOR2X1TS U5978 ( .A(n9949), .B(n12401), .Y(n6255) );
  OAI211X1TS U5975 ( .A0(n12425), .A1(n10166), .B0(n6519), .C0(n5716), .Y(
        n6515) );
  AOI22X1TS U5973 ( .A0(n12240), .A1(n11699), .B0(n11014), .B1(n5551), .Y(
        n6517) );
  OAI21X1TS U6601 ( .A0(n11972), .A1(n12272), .B0(n9962), .Y(n6518) );
  OAI211X1TS U5972 ( .A0(n11287), .A1(n12041), .B0(n6517), .C0(n6518), .Y(
        n6516) );
  NOR3X1TS U5971 ( .A(n6514), .B(n6515), .C(n6516), .Y(n5496) );
  NOR2X1TS U6579 ( .A(n11704), .B(n11013), .Y(n5528) );
  OAI22X1TS U5302 ( .A0(n5528), .A1(n10929), .B0(n11300), .B1(n11305), .Y(
        n5498) );
  NOR2X1TS U5301 ( .A(n10169), .B(n11294), .Y(n5389) );
  OAI22X1TS U5300 ( .A0(n5523), .A1(n10165), .B0(n5389), .B1(n11289), .Y(n5499) );
  NOR2X1TS U6607 ( .A(n10470), .B(n11306), .Y(n5520) );
  NOR2X1TS U5299 ( .A(n10925), .B(n9706), .Y(n5521) );
  OAI211X1TS U5297 ( .A0(n9303), .A1(n10924), .B0(n5518), .C0(n5519), .Y(n5500) );
  NOR2X1TS U6585 ( .A(n9706), .B(n9774), .Y(n5910) );
  NOR4BX1TS U5486 ( .AN(n5909), .B(n5910), .C(n5911), .D(n5912), .Y(n5502) );
  NOR2X1TS U5626 ( .A(n10918), .B(n11389), .Y(n5509) );
  INVX2TS U5289 ( .A(n9170), .Y(n5190) );
  NOR2X1TS U6448 ( .A(n11263), .B(n11205), .Y(n5878) );
  NOR2X1TS U6381 ( .A(n11383), .B(n11239), .Y(n5879) );
  NOR2X1TS U6461 ( .A(n6202), .B(n6779), .Y(n6229) );
  NOR2X1TS U5686 ( .A(n9334), .B(n12383), .Y(n5880) );
  NOR4BX1TS U5467 ( .AN(n5877), .B(n5878), .C(n5879), .D(n5880), .Y(n5868) );
  NOR2X1TS U6517 ( .A(n9836), .B(n9326), .Y(n6784) );
  OAI22X1TS U5466 ( .A0(n9330), .A1(n12415), .B0(n9335), .B1(n10531), .Y(n5873) );
  INVX2TS U6504 ( .A(n9436), .Y(n5861) );
  OAI32X1TS U5465 ( .A0(n5873), .A1(n11276), .A2(n11210), .B0(n11686), .B1(
        n5873), .Y(n5869) );
  NOR2X1TS U5464 ( .A(n10436), .B(n12418), .Y(n5686) );
  NOR2X1TS U6489 ( .A(n12511), .B(n10884), .Y(n5872) );
  OAI22X1TS U5463 ( .A0(n5872), .A1(n10526), .B0(n10857), .B1(n11384), .Y(
        n5871) );
  INVX2TS U6392 ( .A(n12502), .Y(n6087) );
  AOI22X1TS U5868 ( .A0(n10862), .A1(n6217), .B0(n10457), .B1(n11680), .Y(
        n6415) );
  NOR2X1TS U6449 ( .A(n9330), .B(n10427), .Y(n6417) );
  NOR2X1TS U6411 ( .A(n10157), .B(n10431), .Y(n6418) );
  OAI211X1TS U5866 ( .A0(n10213), .A1(n10436), .B0(n6415), .C0(n6416), .Y(
        n6414) );
  OAI211X1TS U5863 ( .A0(n10890), .A1(n10427), .B0(n6412), .C0(n6057), .Y(
        n5467) );
  NOR2X1TS U5895 ( .A(n10529), .B(n11240), .Y(n6436) );
  NOR2X1TS U5894 ( .A(n9330), .B(n11383), .Y(n6216) );
  OAI211X1TS U5886 ( .A0(n6433), .A1(n10432), .B0(n6434), .C0(n6435), .Y(n5468) );
  NOR2X1TS U6446 ( .A(n9945), .B(n12415), .Y(n5487) );
  NOR2X1TS U5849 ( .A(n10161), .B(n11681), .Y(n5457) );
  AOI22X1TS U5283 ( .A0(n11270), .A1(n5480), .B0(n12263), .B1(n5485), .Y(n5471) );
  AOI22X1TS U5282 ( .A0(n11688), .A1(n5480), .B0(n9957), .B1(n9297), .Y(n5472)
         );
  NOR2X1TS U6415 ( .A(n11245), .B(n12033), .Y(n6068) );
  NOR2X1TS U6391 ( .A(n6068), .B(n6087), .Y(n5475) );
  NOR2X1TS U6426 ( .A(n12581), .B(n12264), .Y(n5477) );
  NOR2X1TS U5712 ( .A(n10422), .B(n6229), .Y(n5348) );
  AOI211X1TS U5280 ( .A0(n12219), .A1(n5474), .B0(n5475), .C0(n5476), .Y(n5473) );
  NOR2X1TS U6425 ( .A(n12265), .B(n10458), .Y(n6070) );
  NOR2X1TS U6398 ( .A(n10581), .B(n11233), .Y(n6432) );
  OAI32X1TS U5881 ( .A0(n6427), .A1(n11687), .A2(n11975), .B0(n10863), .B1(
        n6427), .Y(n5429) );
  OAI211X1TS U5904 ( .A0(n11204), .A1(n11258), .B0(n6449), .C0(n6450), .Y(
        n6442) );
  NOR2X1TS U5903 ( .A(n9945), .B(n12386), .Y(n6215) );
  OAI211X1TS U5900 ( .A0(n12417), .A1(n10158), .B0(n6447), .C0(n5691), .Y(
        n6443) );
  AOI22X1TS U5898 ( .A0(n12217), .A1(n11681), .B0(n11000), .B1(n5485), .Y(
        n6445) );
  OAI21X1TS U6406 ( .A0(n11975), .A1(n12263), .B0(n9958), .Y(n6446) );
  OAI211X1TS U5897 ( .A0(n11239), .A1(n12025), .B0(n6445), .C0(n6446), .Y(
        n6444) );
  NOR3X1TS U5896 ( .A(n6442), .B(n6443), .C(n6444), .Y(n5430) );
  NOR2X1TS U6384 ( .A(n11686), .B(n11001), .Y(n5462) );
  OAI22X1TS U5277 ( .A0(n5462), .A1(n10903), .B0(n11252), .B1(n11258), .Y(
        n5432) );
  NOR2X1TS U5276 ( .A(n10161), .B(n11246), .Y(n5350) );
  OAI22X1TS U5275 ( .A0(n5457), .A1(n10157), .B0(n5350), .B1(n11241), .Y(n5433) );
  NOR2X1TS U6412 ( .A(n10461), .B(n11258), .Y(n5454) );
  NOR2X1TS U5274 ( .A(n10898), .B(n9702), .Y(n5455) );
  OAI211X1TS U5272 ( .A0(n9293), .A1(n10897), .B0(n5452), .C0(n5453), .Y(n5434) );
  NOR2X1TS U6390 ( .A(n9702), .B(n9770), .Y(n5854) );
  OAI22X1TS U5458 ( .A0(n11359), .A1(n10891), .B0(n10505), .B1(n10209), .Y(
        n5855) );
  NOR4BX1TS U5453 ( .AN(n5853), .B(n5854), .C(n5855), .D(n5856), .Y(n5436) );
  NOR2X1TS U5598 ( .A(n10890), .B(n11383), .Y(n5443) );
  INVX2TS U5264 ( .A(n9145), .Y(n5123) );
  NOR2X1TS U6939 ( .A(n6918), .B(n10721), .Y(n6901) );
  NOR2X1TS U6908 ( .A(sa01[6]), .B(n6318), .Y(n6904) );
  NOR2X1TS U6913 ( .A(n9452), .B(sa01[4]), .Y(n6905) );
  AOI22X1TS U6158 ( .A0(n5745), .A1(n12543), .B0(n11724), .B1(n11355), .Y(
        n6641) );
  INVX2TS U6918 ( .A(n6338), .Y(n6911) );
  INVX2TS U6879 ( .A(n6351), .Y(n5753) );
  INVX2TS U6912 ( .A(n6317), .Y(n6674) );
  INVX2TS U6916 ( .A(n6897), .Y(n6319) );
  NOR2X1TS U6904 ( .A(n10974), .B(n9782), .Y(n6675) );
  AOI22X1TS U6155 ( .A0(n11997), .A1(n12534), .B0(n10946), .B1(n12434), .Y(
        n6668) );
  AOI22X1TS U6152 ( .A0(n12062), .A1(n12431), .B0(n9978), .B1(n6289), .Y(n6669) );
  INVX2TS U6892 ( .A(n9397), .Y(n6639) );
  AOI21X1TS U6149 ( .A0(n10964), .A1(n6633), .B0(n6671), .Y(n6670) );
  NOR2X1TS U6824 ( .A(n11999), .B(n12542), .Y(n5759) );
  OAI22X1TS U6147 ( .A0(n5759), .A1(n11735), .B0(n11746), .B1(n10517), .Y(
        n6666) );
  AOI211X1TS U6146 ( .A0(n12294), .A1(n10177), .B0(n6357), .C0(n6666), .Y(
        n6643) );
  NOR2X1TS U6143 ( .A(n10233), .B(n10488), .Y(n6299) );
  AOI211X1TS U6142 ( .A0(n10249), .A1(n10181), .B0(n6665), .C0(n6299), .Y(
        n6663) );
  OAI211X1TS U6141 ( .A0(n11746), .A1(n10234), .B0(n6663), .C0(n6664), .Y(
        n6662) );
  NOR2X1TS U6139 ( .A(n6320), .B(n11983), .Y(n6279) );
  AOI221X1TS U6138 ( .A0(n12545), .A1(n5954), .B0(n10238), .B1(n12298), .C0(
        n6279), .Y(n6661) );
  OAI211X1TS U6137 ( .A0(n12020), .A1(n9403), .B0(n6660), .C0(n6661), .Y(n6326) );
  NOR2X1TS U6127 ( .A(n10545), .B(n12537), .Y(n5589) );
  NOR2X1TS U6830 ( .A(n12544), .B(n11354), .Y(n6631) );
  INVX2TS U6829 ( .A(n6631), .Y(n6286) );
  AOI22X1TS U6125 ( .A0(n10194), .A1(n5988), .B0(n5959), .B1(n6286), .Y(n6650)
         );
  AOI22X1TS U6122 ( .A0(n12280), .A1(n6649), .B0(n11353), .B1(n5962), .Y(n6647) );
  NOR2X1TS U6115 ( .A(n9973), .B(n12300), .Y(n5597) );
  AOI31X1TS U6114 ( .A0(n5597), .A1(n9981), .A2(n12287), .B0(n12005), .Y(n6636) );
  OAI211X1TS U6110 ( .A0(n6311), .A1(n11753), .B0(n6634), .C0(n6635), .Y(n6601) );
  NOR2X1TS U6109 ( .A(n11347), .B(n12543), .Y(n5674) );
  NOR2X1TS U6840 ( .A(n10483), .B(n9403), .Y(n6623) );
  AOI22X1TS U6106 ( .A0(n11718), .A1(n12299), .B0(n10550), .B1(n11330), .Y(
        n6625) );
  OAI21X1TS U6105 ( .A0(n10968), .A1(n10181), .B0(n12056), .Y(n6626) );
  AOI211X1TS U6101 ( .A0(n10576), .A1(n12536), .B0(n6628), .C0(n6629), .Y(
        n6627) );
  AOI211X1TS U6099 ( .A0(n12431), .A1(n12056), .B0(n6623), .C0(n6330), .Y(
        n6622) );
  OAI211X1TS U6098 ( .A0(n5674), .A1(n12021), .B0(n6621), .C0(n6622), .Y(n6602) );
  AOI22X1TS U6091 ( .A0(n10576), .A1(n5959), .B0(n12292), .B1(n6295), .Y(n6606) );
  OAI21X1TS U6089 ( .A0(n11717), .A1(n10202), .B0(n10963), .Y(n6613) );
  OAI211X1TS U6088 ( .A0(n11983), .A1(n12006), .B0(n5970), .C0(n6613), .Y(
        n6607) );
  OAI21X1TS U6086 ( .A0(n11348), .A1(n10182), .B0(n5760), .Y(n6612) );
  NOR4BX1TS U6080 ( .AN(n6606), .B(n6607), .C(n6608), .D(n6609), .Y(n5765) );
  OAI21X1TS U6079 ( .A0(n5599), .A1(n12299), .B0(n12292), .Y(n6604) );
  AOI22X1TS U6078 ( .A0(n11349), .A1(n10479), .B0(n10202), .B1(n10250), .Y(
        n6605) );
  NOR2X1TS U6347 ( .A(n6049), .B(sa30[6]), .Y(n6542) );
  NOR2X1TS U6345 ( .A(n9429), .B(n10327), .Y(n6737) );
  NOR2X1TS U6338 ( .A(n9819), .B(n10715), .Y(n6720) );
  AOI22X1TS U6335 ( .A0(n10840), .A1(n9993), .B0(n11397), .B1(n11337), .Y(
        n6703) );
  NOR2X1TS U6331 ( .A(n10043), .B(n9812), .Y(n5625) );
  NOR2X1TS U6321 ( .A(n10043), .B(n6049), .Y(n6738) );
  NOR2X1TS U6315 ( .A(n10190), .B(n9762), .Y(n6532) );
  INVX2TS U6303 ( .A(n9747), .Y(n6702) );
  AOI22X1TS U6297 ( .A0(n11342), .A1(n6699), .B0(n11697), .B1(n11337), .Y(
        n6735) );
  NOR2X1TS U6290 ( .A(n10818), .B(n12210), .Y(n6554) );
  NOR2X1TS U6287 ( .A(n10413), .B(n10522), .Y(n6572) );
  AOI211X1TS U6286 ( .A0(n11670), .A1(n6027), .B0(n6554), .C0(n6572), .Y(n6736) );
  OAI22X1TS U6277 ( .A0(n5632), .A1(n12497), .B0(n12442), .B1(n10185), .Y(
        n6731) );
  AOI211X1TS U6276 ( .A0(n10245), .A1(n11981), .B0(n6168), .C0(n6731), .Y(
        n6705) );
  AOI22X1TS U6274 ( .A0(n11227), .A1(n11679), .B0(n11395), .B1(n11341), .Y(
        n6725) );
  NOR2X1TS U6266 ( .A(n10989), .B(n10847), .Y(n6030) );
  AOI211X1TS U6265 ( .A0(n10554), .A1(n10497), .B0(n6729), .C0(n6030), .Y(
        n6726) );
  OAI32X1TS U6254 ( .A0(n6723), .A1(n9376), .A2(n12448), .B0(n11685), .B1(
        n6723), .Y(n6722) );
  OAI211X1TS U6251 ( .A0(n12441), .A1(n10990), .B0(n6722), .C0(n6560), .Y(
        n6142) );
  NOR2X1TS U6248 ( .A(n9969), .B(n10242), .Y(n5413) );
  INVX2TS U6247 ( .A(n5413), .Y(n6162) );
  AOI22X1TS U6246 ( .A0(n11685), .A1(n10952), .B0(n11336), .B1(n6162), .Y(
        n6711) );
  NOR2X1TS U6244 ( .A(n12203), .B(n10846), .Y(n6531) );
  OAI32X1TS U6242 ( .A0(n6531), .A1(n9953), .A2(n11695), .B0(n11377), .B1(
        n6531), .Y(n6712) );
  OAI21X1TS U6237 ( .A0(n10841), .A1(n10497), .B0(n11396), .Y(n6718) );
  AOI32X1TS U6236 ( .A0(n10984), .A1(n6718), .A2(n9758), .B0(n12205), .B1(
        n6718), .Y(n6716) );
  AOI211X1TS U6233 ( .A0(n10492), .A1(n6715), .B0(n6716), .C0(n6717), .Y(n6713) );
  NOR2X1TS U6229 ( .A(n11397), .B(n9994), .Y(n6028) );
  AOI22X1TS U6224 ( .A0(n11378), .A1(n6584), .B0(n10241), .B1(n5808), .Y(n6710) );
  AOI22X1TS U6219 ( .A0(n11683), .A1(n6580), .B0(n9994), .B1(n5785), .Y(n6709)
         );
  NOR2X1TS U6210 ( .A(n11379), .B(n11229), .Y(n5315) );
  NOR2X1TS U6202 ( .A(n11676), .B(n9989), .Y(n6544) );
  OAI22X1TS U6201 ( .A0(n6028), .A1(n10154), .B0(n6544), .B1(n10989), .Y(n6691) );
  OAI22X1TS U6200 ( .A0(n11403), .A1(n11977), .B0(n10959), .B1(n10830), .Y(
        n6692) );
  AOI21X1TS U6199 ( .A0(n12442), .A1(n11691), .B0(n10189), .Y(n6693) );
  NOR2X1TS U6198 ( .A(n10150), .B(n10818), .Y(n6570) );
  NOR2X1TS U6197 ( .A(n10847), .B(n10979), .Y(n6020) );
  OAI211X1TS U6194 ( .A0(n10984), .A1(n12198), .B0(n6695), .C0(n6696), .Y(
        n6694) );
  NOR2X1TS U6191 ( .A(n10417), .B(n9759), .Y(n6578) );
  NOR2X1TS U6190 ( .A(n11396), .B(n11674), .Y(n5414) );
  NOR2X1TS U6186 ( .A(n10819), .B(n6010), .Y(n6591) );
  NOR2X1TS U6184 ( .A(n10416), .B(n10412), .Y(n6575) );
  NOR2X1TS U6183 ( .A(n10991), .B(n10825), .Y(n6587) );
  AOI211X1TS U6182 ( .A0(n10491), .A1(n6581), .B0(n6575), .C0(n6587), .Y(n6688) );
  OAI211X1TS U6180 ( .A0(n9766), .A1(n10153), .B0(n6688), .C0(n6029), .Y(n6687) );
  AOI211X1TS U6179 ( .A0(n10142), .A1(n9997), .B0(n6591), .C0(n6687), .Y(n6163) );
  NOR2X1TS U6178 ( .A(n12450), .B(n10834), .Y(n6014) );
  OAI22X1TS U6177 ( .A0(n6014), .A1(n9767), .B0(n11402), .B1(n10413), .Y(n6681) );
  OAI21X1TS U6171 ( .A0(n11207), .A1(n9970), .B0(n11343), .Y(n6686) );
  OAI21X1TS U6168 ( .A0(n10554), .A1(n11675), .B0(n10836), .Y(n6685) );
  OAI211X1TS U6166 ( .A0(n11977), .A1(n10501), .B0(n6685), .C0(n5422), .Y(
        n6684) );
  OAI22X1TS U5245 ( .A0(n5387), .A1(n10452), .B0(n5389), .B1(n9949), .Y(n5386)
         );
  AOI211X1TS U5244 ( .A0(n12590), .A1(n10440), .B0(n5385), .C0(n5386), .Y(
        n5383) );
  OAI211X1TS U5243 ( .A0(n5380), .A1(n12401), .B0(n5382), .C0(n5383), .Y(n5357) );
  AOI22X1TS U5242 ( .A0(n12242), .A1(n10880), .B0(n12248), .B1(n5379), .Y(
        n5374) );
  OAI211X1TS U5241 ( .A0(n5506), .A1(n10449), .B0(n5374), .C0(n5375), .Y(n5358) );
  OAI22X1TS U5925 ( .A0(n5543), .A1(n11366), .B0(n6467), .B1(n10540), .Y(n6461) );
  OAI22X1TS U5923 ( .A0(n5523), .A1(n11300), .B0(n9367), .B1(n12425), .Y(n6462) );
  AOI22X1TS U5920 ( .A0(n11705), .A1(n9734), .B0(n10912), .B1(n12521), .Y(
        n6465) );
  AOI32X1TS U5919 ( .A0(n6465), .A1(n11215), .A2(n11301), .B0(n10222), .B1(
        n6465), .Y(n6464) );
  NOR2X1TS U5935 ( .A(n10512), .B(n10444), .Y(n6249) );
  NOR2X1TS U6722 ( .A(n5558), .B(n10572), .Y(n6478) );
  OAI21X1TS U5934 ( .A0(n11705), .A1(n11414), .B0(n12249), .Y(n6479) );
  AOI22X1TS U5933 ( .A0(n10935), .A1(n10914), .B0(n11704), .B1(n11008), .Y(
        n6480) );
  AOI211X1TS U5931 ( .A0(n11282), .A1(n10878), .B0(n6249), .C0(n6477), .Y(
        n5361) );
  NOR2X1TS U6640 ( .A(n10222), .B(n11288), .Y(n5889) );
  OAI22X1TS U5480 ( .A0(n5899), .A1(n9950), .B0(n11299), .B1(n11391), .Y(n5890) );
  AOI21X1TS U5477 ( .A0(n11299), .A1(n10452), .B0(n10924), .Y(n5896) );
  OAI32X1TS U5476 ( .A0(n5896), .A1(n11295), .A2(n12249), .B0(n10936), .B1(
        n5896), .Y(n5893) );
  INVX2TS U5203 ( .A(n9279), .Y(n1582) );
  AOI22X1TS U7435 ( .A0(n11914), .A1(n7698), .B0(n12142), .B1(n11138), .Y(
        n7817) );
  AOI22X1TS U7434 ( .A0(n12191), .A1(n9869), .B0(n11861), .B1(n12618), .Y(
        n7818) );
  AOI22X1TS U7433 ( .A0(n12370), .A1(n7825), .B0(n12364), .B1(n7826), .Y(n7819) );
  OAI21X1TS U7432 ( .A0(n12357), .A1(n10661), .B0(n7823), .Y(n7822) );
  AOI211X1TS U7431 ( .A0(n11593), .A1(n12363), .B0(n7821), .C0(n7822), .Y(
        n7820) );
  OAI22X1TS U7356 ( .A0(n11904), .A1(n10707), .B0(n10073), .B1(n9858), .Y(
        n7697) );
  OAI211X1TS U7449 ( .A0(n7854), .A1(n11528), .B0(n7855), .C0(n7856), .Y(n7853) );
  NOR3X1TS U7448 ( .A(n7851), .B(n7852), .C(n7853), .Y(n7677) );
  OAI22X1TS U7330 ( .A0(n7667), .A1(n11598), .B0(n7494), .B1(n9846), .Y(n7636)
         );
  AOI22X1TS U7328 ( .A0(n12632), .A1(n7663), .B0(n12185), .B1(n7664), .Y(n7660) );
  AOI211X1TS U7321 ( .A0(n11916), .A1(n12349), .B0(n7646), .C0(n7647), .Y(
        n7642) );
  INVX2TS U7317 ( .A(n9224), .Y(n6976) );
  AOI22X1TS U7225 ( .A0(n6976), .A1(n9480), .B0(n9478), .B1(n9224), .Y(n7344)
         );
  OAI22X1TS U7188 ( .A0(n7367), .A1(n11806), .B0(n11112), .B1(n7230), .Y(n7362) );
  OAI22X1TS U7187 ( .A0(n9830), .A1(n10266), .B0(n7365), .B1(n11874), .Y(n7363) );
  AOI22X1TS U7480 ( .A0(n11565), .A1(n10018), .B0(n10253), .B1(n10324), .Y(
        n7874) );
  AOI211X1TS U7473 ( .A0(n11445), .A1(n7878), .B0(n7524), .C0(n7879), .Y(n7876) );
  AOI22X1TS U7184 ( .A0(n11534), .A1(n11451), .B0(n11038), .B1(n10254), .Y(
        n7355) );
  OAI22X1TS U7175 ( .A0(n7340), .A1(n12734), .B0(n12682), .B1(n7341), .Y(N113)
         );
  OAI22X1TS U3352 ( .A0(n3550), .A1(n10480), .B0(n3552), .B1(n9915), .Y(n3549)
         );
  AOI211X1TS U3351 ( .A0(n12586), .A1(n10494), .B0(n3548), .C0(n3549), .Y(
        n3546) );
  OAI211X1TS U3350 ( .A0(n3543), .A1(n12445), .B0(n3545), .C0(n3546), .Y(n3520) );
  AOI22X1TS U3349 ( .A0(n12269), .A1(n10907), .B0(n12260), .B1(n3542), .Y(
        n3537) );
  OAI211X1TS U3348 ( .A0(n3685), .A1(n10486), .B0(n3537), .C0(n3538), .Y(n3521) );
  OAI22X1TS U3967 ( .A0(n3722), .A1(n11262), .B0(n4595), .B1(n10392), .Y(n4589) );
  OAI22X1TS U3965 ( .A0(n3702), .A1(n11351), .B0(n9153), .B1(n12405), .Y(n4590) );
  AOI22X1TS U3962 ( .A0(n11745), .A1(n9646), .B0(n10854), .B1(n12525), .Y(
        n4593) );
  AOI32X1TS U3961 ( .A0(n4593), .A1(n11410), .A2(n11351), .B0(n10110), .B1(
        n4593), .Y(n4592) );
  NOR2X1TS U3977 ( .A(n10424), .B(n10489), .Y(n4406) );
  NOR2X1TS U4644 ( .A(n3737), .B(n10377), .Y(n4606) );
  OAI21X1TS U3976 ( .A0(n11744), .A1(n11230), .B0(n12261), .Y(n4607) );
  AOI22X1TS U3975 ( .A0(n10833), .A1(n10856), .B0(n11743), .B1(n10762), .Y(
        n4608) );
  AOI211X1TS U3973 ( .A0(n11369), .A1(n10907), .B0(n4406), .C0(n4605), .Y(
        n3524) );
  NOR2X1TS U4562 ( .A(n10109), .B(n11362), .Y(n4033) );
  OAI22X1TS U3564 ( .A0(n4043), .A1(n9916), .B0(n11350), .B1(n11244), .Y(n4034) );
  AOI21X1TS U3561 ( .A0(n11350), .A1(n10480), .B0(n10844), .Y(n4040) );
  OAI32X1TS U3560 ( .A0(n4040), .A1(n11356), .A2(n12262), .B0(n10832), .B1(
        n4040), .Y(n4037) );
  AOI22X1TS U3923 ( .A0(n11213), .A1(n12032), .B0(n10806), .B1(n4324), .Y(
        n4541) );
  NOR2X1TS U3921 ( .A(n10866), .B(n10456), .Y(n4327) );
  AOI211X1TS U3920 ( .A0(n10410), .A1(n9679), .B0(n4543), .C0(n4327), .Y(n4542) );
  OAI211X1TS U3919 ( .A0(n10790), .A1(n9676), .B0(n4541), .C0(n4542), .Y(n4540) );
  OAI22X1TS U3515 ( .A0(n11762), .A1(n12379), .B0(n12207), .B1(n11715), .Y(
        n3942) );
  OAI22X1TS U3514 ( .A0(n3953), .A1(n12540), .B0(n3954), .B1(n12412), .Y(n3943) );
  NOR2X1TS U4921 ( .A(n10771), .B(n9921), .Y(n3951) );
  NOR2X1TS U4886 ( .A(n10111), .B(n9675), .Y(n3952) );
  AOI211X1TS U3513 ( .A0(n10410), .A1(n3911), .B0(n3951), .C0(n3952), .Y(n3945) );
  OAI22X1TS U3512 ( .A0(n10112), .A1(n12022), .B0(n9650), .B1(n12413), .Y(
        n3948) );
  OAI211X1TS U3510 ( .A0(n12568), .A1(n12539), .B0(n3945), .C0(n3946), .Y(
        n3944) );
  NOR3X1TS U3509 ( .A(n3942), .B(n3943), .C(n3944), .Y(n3632) );
  OAI22X1TS U3392 ( .A0(n10144), .A1(n3663), .B0(n11757), .B1(n12532), .Y(
        n3655) );
  OAI22X1TS U3391 ( .A0(n11763), .A1(n12541), .B0(n4480), .B1(n10455), .Y(
        n3656) );
  AOI22X1TS U4926 ( .A0(n10116), .A1(n9686), .B0(n4841), .B1(n9190), .Y(n3641)
         );
  OAI211X1TS U3384 ( .A0(n3639), .A1(n11774), .B0(n3641), .C0(n3642), .Y(n3638) );
  OAI22X1TS U5234 ( .A0(n5348), .A1(n10435), .B0(n5350), .B1(n9945), .Y(n5347)
         );
  AOI211X1TS U5233 ( .A0(n12581), .A1(n10422), .B0(n5346), .C0(n5347), .Y(
        n5344) );
  OAI211X1TS U5232 ( .A0(n5341), .A1(n12385), .B0(n5343), .C0(n5344), .Y(n5318) );
  AOI22X1TS U5231 ( .A0(n12219), .A1(n10863), .B0(n12225), .B1(n5340), .Y(
        n5335) );
  OAI211X1TS U5230 ( .A0(n5440), .A1(n10432), .B0(n5335), .C0(n5336), .Y(n5319) );
  OAI22X1TS U5850 ( .A0(n5477), .A1(n11360), .B0(n6395), .B1(n10531), .Y(n6389) );
  OAI22X1TS U5848 ( .A0(n5457), .A1(n11252), .B0(n9359), .B1(n12417), .Y(n6390) );
  AOI22X1TS U5845 ( .A0(n11687), .A1(n9730), .B0(n10886), .B1(n12504), .Y(
        n6393) );
  NOR2X1TS U5860 ( .A(n10506), .B(n10427), .Y(n6209) );
  NOR2X1TS U6527 ( .A(n5492), .B(n10567), .Y(n6406) );
  OAI21X1TS U5859 ( .A0(n11687), .A1(n11407), .B0(n12225), .Y(n6407) );
  AOI22X1TS U5858 ( .A0(n5874), .A1(n10885), .B0(n11686), .B1(n10996), .Y(
        n6408) );
  AOI211X1TS U5856 ( .A0(n11234), .A1(n10862), .B0(n6209), .C0(n6405), .Y(
        n5322) );
  NOR2X1TS U6445 ( .A(n10214), .B(n11241), .Y(n5833) );
  OAI22X1TS U5447 ( .A0(n5843), .A1(n9946), .B0(n11251), .B1(n11384), .Y(n5834) );
  AOI21X1TS U5444 ( .A0(n11251), .A1(n10435), .B0(n10897), .Y(n5840) );
  OAI32X1TS U5443 ( .A0(n5840), .A1(n11246), .A2(n12226), .B0(n10909), .B1(
        n5840), .Y(n5837) );
  OAI22X1TS U5403 ( .A0(n11729), .A1(n10518), .B0(n11371), .B1(n11754), .Y(
        n5747) );
  OAI22X1TS U5402 ( .A0(n5759), .A1(n12286), .B0(n11730), .B1(n10473), .Y(
        n5748) );
  NOR2X1TS U6809 ( .A(n9727), .B(n9781), .Y(n5757) );
  NOR2X1TS U6770 ( .A(n10197), .B(n10226), .Y(n5758) );
  AOI211X1TS U5401 ( .A0(n10201), .A1(n5670), .B0(n5757), .C0(n5758), .Y(n5751) );
  OAI211X1TS U5398 ( .A0(n11747), .A1(n12285), .B0(n5751), .C0(n5752), .Y(
        n5749) );
  NOR3X1TS U5397 ( .A(n5747), .B(n5748), .C(n5749), .Y(n5561) );
  AOI211X1TS U5801 ( .A0(n10964), .A1(n10193), .B0(n6346), .C0(n6347), .Y(
        n6344) );
  INVX2TS U6859 ( .A(n12278), .Y(n6334) );
  AOI32X1TS U5323 ( .A0(n5597), .A1(n5598), .A2(n10484), .B0(n5743), .B1(n5598), .Y(n5587) );
  AOI22X1TS U6816 ( .A0(n10193), .A1(n10941), .B0(n9974), .B1(n10237), .Y(
        n5591) );
  AOI211X1TS U5320 ( .A0(n10947), .A1(n5586), .B0(n5587), .C0(n5588), .Y(n5565) );
  AOI22X1TS U5319 ( .A0(n12545), .A1(n10479), .B0(n10182), .B1(n10942), .Y(
        n5566) );
  AOI22X1TS U5318 ( .A0(n12433), .A1(n10178), .B0(n11330), .B1(n12537), .Y(
        n5567) );
  NOR2X1TS U5755 ( .A(n10198), .B(n5585), .Y(n5569) );
  NOR2X1TS U5773 ( .A(n9982), .B(n9778), .Y(n5570) );
  OAI21X1TS U5818 ( .A0(n11347), .A1(n10238), .B0(n9977), .Y(n6367) );
  NOR2X1TS U6844 ( .A(n11998), .B(n11354), .Y(n5973) );
  AOI22X1TS U5817 ( .A0(n12056), .A1(n9352), .B0(n12535), .B1(n6372), .Y(n6368) );
  NOR2X1TS U6792 ( .A(n9726), .B(n9388), .Y(n6370) );
  AOI211X1TS U5815 ( .A0(n11716), .A1(n10940), .B0(n6370), .C0(n6371), .Y(
        n6369) );
  NOR4BX1TS U5314 ( .AN(n5561), .B(n5562), .C(n5563), .D(n5564), .Y(n5122) );
  INVX2TS U5222 ( .A(n5122), .Y(n1778) );
  NOR2X1TS U5651 ( .A(n9965), .B(n10206), .Y(n5419) );
  NOR2X1TS U5650 ( .A(n10979), .B(n9767), .Y(n6016) );
  AOI211X1TS U5649 ( .A0(n10245), .A1(n9970), .B0(n5419), .C0(n6016), .Y(n6156) );
  AOI31X1TS U5648 ( .A0(n12440), .A1(n9762), .A2(n11673), .B0(n12497), .Y(
        n6158) );
  AOI211X1TS U5645 ( .A0(n10835), .A1(n11396), .B0(n6158), .C0(n6159), .Y(
        n6157) );
  NOR2X1TS U6030 ( .A(n10522), .B(n9763), .Y(n5618) );
  OAI22X1TS U5344 ( .A0(n5632), .A1(n12198), .B0(n11976), .B1(n10959), .Y(
        n5619) );
  OAI22X1TS U5343 ( .A0(n5411), .A1(n12211), .B0(n9966), .B1(n11673), .Y(n5620) );
  AOI22X1TS U5342 ( .A0(n10492), .A1(n10497), .B0(n11695), .B1(n11669), .Y(
        n5623) );
  OAI22X1TS U5341 ( .A0(n12205), .A1(n11671), .B0(n11978), .B1(n10186), .Y(
        n5627) );
  AOI32X1TS U5220 ( .A0(n5313), .A1(n6024), .A2(n5315), .B0(n10846), .B1(n5313), .Y(n5303) );
  AOI22X1TS U6049 ( .A0(n9376), .A1(n10242), .B0(n10492), .B1(n11227), .Y(
        n5308) );
  OAI211X1TS U5218 ( .A0(n5305), .A1(n12209), .B0(n5307), .C0(n5308), .Y(n5304) );
  AOI211X1TS U5217 ( .A0(n10836), .A1(n9283), .B0(n5303), .C0(n5304), .Y(n5278) );
  OAI22X1TS U5216 ( .A0(n12496), .A1(n11691), .B0(n12203), .B1(n10150), .Y(
        n5281) );
  OAI22X1TS U5215 ( .A0(n10826), .A1(n12197), .B0(n10829), .B1(n9942), .Y(
        n5282) );
  NOR2X1TS U5544 ( .A(n11671), .B(n10186), .Y(n5292) );
  AOI221X1TS U5214 ( .A0(n6161), .A1(n10141), .B0(n11697), .B1(n10146), .C0(
        n5292), .Y(n5286) );
  INVX2TS U5664 ( .A(n9312), .Y(n5784) );
  INVX2TS U5210 ( .A(n9203), .Y(n5132) );
  INVX2TS U5208 ( .A(n5191), .Y(n5192) );
  AOI211X1TS U7098 ( .A0(n11449), .A1(n11456), .B0(n7142), .C0(n7143), .Y(
        n7139) );
  NOR4BX1TS U7092 ( .AN(n7115), .B(n7116), .C(n7117), .D(n7118), .Y(n7102) );
  AOI211X1TS U7089 ( .A0(n10254), .A1(n10258), .B0(n7107), .C0(n7108), .Y(
        n7103) );
  NOR4X1TS U7087 ( .A(n7097), .B(n7098), .C(n7099), .D(n7100), .Y(n1602) );
  INVX2TS U7086 ( .A(n1602), .Y(n1604) );
  OAI22X1TS U7012 ( .A0(n1604), .A1(n1562), .B0(n1563), .B1(n1602), .Y(n1278)
         );
  OAI22X1TS U8771 ( .A0(n11820), .A1(n11777), .B0(n9467), .B1(n11467), .Y(
        n8672) );
  OAI22X1TS U8743 ( .A0(n11604), .A1(n11836), .B0(n11832), .B1(n11425), .Y(
        n8674) );
  AOI21X1TS U8738 ( .A0(n11421), .A1(n10601), .B0(n12149), .Y(n8675) );
  AOI32X1TS U8734 ( .A0(n7937), .A1(n8669), .A2(n12328), .B0(n11766), .B1(
        n8669), .Y(n7907) );
  AOI22X1TS U8631 ( .A0(n11880), .A1(n11053), .B0(n11825), .B1(n11048), .Y(
        n8625) );
  AOI22X1TS U8627 ( .A0(n11826), .A1(n7789), .B0(n10290), .B1(n7394), .Y(n8627) );
  AOI22X1TS U8615 ( .A0(n11879), .A1(n7215), .B0(n11940), .B1(n7789), .Y(n8617) );
  AOI211X1TS U8613 ( .A0(n11784), .A1(n8158), .B0(n8615), .C0(n8616), .Y(n8614) );
  OAI22X1TS U7006 ( .A0(n6992), .A1(n12739), .B0(n12683), .B1(n6993), .Y(N132)
         );
  NOR2X1TS U6519 ( .A(n12218), .B(n10851), .Y(n6195) );
  AOI22X1TS U6498 ( .A0(n11245), .A1(n11687), .B0(n12227), .B1(n11235), .Y(
        n6796) );
  NOR2X1TS U6491 ( .A(n10213), .B(n10507), .Y(n5828) );
  AOI211X1TS U6470 ( .A0(n12224), .A1(n10457), .B0(n6789), .C0(n6790), .Y(
        n6788) );
  AOI211X1TS U6467 ( .A0(n12583), .A1(n10162), .B0(n5828), .C0(n6787), .Y(
        n5689) );
  AOI21X1TS U6459 ( .A0(n10158), .A1(n9702), .B0(n12383), .Y(n6422) );
  AOI22X1TS U6452 ( .A0(n11234), .A1(n12035), .B0(n11409), .B1(n11680), .Y(
        n6783) );
  OAI21X1TS U6451 ( .A0(n11264), .A1(n11240), .B0(n6783), .Y(n6782) );
  OAI22X1TS U6436 ( .A0(n10214), .A1(n10526), .B0(n10431), .B1(n10892), .Y(
        n6777) );
  AOI211X1TS U6430 ( .A0(n11235), .A1(n5474), .B0(n6777), .C0(n6778), .Y(n6073) );
  NOR2X1TS U6400 ( .A(n12265), .B(n11001), .Y(n5831) );
  AOI211X1TS U6389 ( .A0(n11408), .A1(n12226), .B0(n5475), .C0(n5854), .Y(
        n6762) );
  OAI22X1TS U6386 ( .A0(n10525), .A1(n10531), .B0(n10436), .B1(n12026), .Y(
        n6757) );
  OAI22X1TS U6383 ( .A0(n6222), .A1(n10568), .B0(n5462), .B1(n11259), .Y(n6758) );
  OAI22X1TS U6380 ( .A0(n11252), .A1(n12027), .B0(n9334), .B1(n11258), .Y(
        n6756) );
  OAI211X1TS U6378 ( .A0(n9292), .A1(n12385), .B0(n6074), .C0(n6075), .Y(n6740) );
  NOR2X1TS U6377 ( .A(n11409), .B(n10457), .Y(n5864) );
  NOR2X1TS U6370 ( .A(n10582), .B(n12582), .Y(n5865) );
  OAI22X1TS U6367 ( .A0(n10567), .A1(n10526), .B0(n10157), .B1(n10904), .Y(
        n6748) );
  OAI22X1TS U6366 ( .A0(n10431), .A1(n11240), .B0(n10505), .B1(n12027), .Y(
        n6749) );
  NOR2X1TS U6365 ( .A(n10422), .B(n9958), .Y(n6388) );
  INVX2TS U6924 ( .A(n6648), .Y(n5989) );
  OAI22X1TS U6895 ( .A0(n6277), .A1(n11734), .B0(n10488), .B1(n11984), .Y(
        n6916) );
  AOI211X1TS U6894 ( .A0(n12536), .A1(n10182), .B0(n6675), .C0(n6916), .Y(
        n5945) );
  NOR2X1TS U6885 ( .A(n11020), .B(n10517), .Y(n6362) );
  NOR2X1TS U6881 ( .A(n10233), .B(n11990), .Y(n5767) );
  AOI211X1TS U6880 ( .A0(n12298), .A1(n12545), .B0(n6362), .C0(n5767), .Y(
        n6907) );
  NOR2X1TS U6871 ( .A(n12294), .B(n10202), .Y(n6315) );
  OAI22X1TS U6869 ( .A0(n6378), .A1(n11729), .B0(n6315), .B1(n10483), .Y(n6913) );
  OAI32X1TS U6865 ( .A0(n6913), .A1(n11722), .A2(n10941), .B0(n10238), .B1(
        n6913), .Y(n6912) );
  OAI211X1TS U6862 ( .A0(n11736), .A1(n10487), .B0(n6912), .C0(n6340), .Y(
        n5950) );
  OAI22X1TS U6853 ( .A0(n6297), .A1(n11752), .B0(n10473), .B1(n10487), .Y(
        n6909) );
  AOI211X1TS U6852 ( .A0(n11718), .A1(n11724), .B0(n5950), .C0(n6909), .Y(
        n6908) );
  OAI211X1TS U6851 ( .A0(n11748), .A1(n11734), .B0(n6907), .C0(n6908), .Y(
        n6857) );
  AOI22X1TS U6837 ( .A0(n12292), .A1(n6649), .B0(n10201), .B1(n6295), .Y(n6903) );
  NOR2X1TS U6827 ( .A(n10550), .B(n10942), .Y(n6374) );
  AOI21X1TS U6820 ( .A0(n10198), .A1(n11989), .B0(n11754), .Y(n6376) );
  AOI211X1TS U6814 ( .A0(n11330), .A1(n6617), .B0(n6376), .C0(n6899), .Y(n6878) );
  NOR2X1TS U6811 ( .A(n10975), .B(n11728), .Y(n5766) );
  AOI22X1TS U6807 ( .A0(n10545), .A1(n12542), .B0(n11722), .B1(n11997), .Y(
        n6898) );
  AOI22X1TS U6805 ( .A0(n10946), .A1(n12292), .B0(n12431), .B1(n12298), .Y(
        n6896) );
  OAI211X1TS U6803 ( .A0(n11747), .A1(n9726), .B0(n6896), .C0(n6364), .Y(n6895) );
  OAI211X1TS U6800 ( .A0(n6892), .A1(n11748), .B0(n6893), .C0(n6664), .Y(n5643) );
  AOI211X1TS U6791 ( .A0(n10193), .A1(n12055), .B0(n6890), .C0(n6370), .Y(
        n6884) );
  OAI211X1TS U6780 ( .A0(n6298), .A1(n12012), .B0(n6884), .C0(n6885), .Y(n5978) );
  AOI22X1TS U6778 ( .A0(n12294), .A1(n10964), .B0(n12432), .B1(n12534), .Y(
        n6883) );
  AOI211X1TS U6771 ( .A0(n12062), .A1(n9353), .B0(n6874), .C0(n6875), .Y(n6272) );
  NOR2X1TS U6765 ( .A(n11353), .B(n11740), .Y(n5746) );
  OAI22X1TS U6764 ( .A0(n5746), .A1(n12013), .B0(n10484), .B1(n10488), .Y(
        n6870) );
  AOI22X1TS U6763 ( .A0(n12054), .A1(n12293), .B0(n11723), .B1(n12433), .Y(
        n6873) );
  OAI22X1TS U6760 ( .A0(n10474), .A1(n12007), .B0(n12021), .B1(n11991), .Y(
        n6864) );
  OAI22X1TS U6758 ( .A0(n11730), .A1(n9722), .B0(n9982), .B1(n10488), .Y(n6865) );
  AOI21X1TS U6757 ( .A0(n12021), .A1(n11735), .B0(n10174), .Y(n6866) );
  AOI22X1TS U6756 ( .A0(n11717), .A1(n6649), .B0(n12063), .B1(n6372), .Y(n6868) );
  NOR2X1TS U6751 ( .A(n11999), .B(n12432), .Y(n5763) );
  NOR2X1TS U6746 ( .A(n10194), .B(n12545), .Y(n5769) );
  AOI22X1TS U6067 ( .A0(n11228), .A1(n9969), .B0(n10555), .B1(n10142), .Y(
        n6593) );
  AOI22X1TS U6064 ( .A0(n11207), .A1(n6580), .B0(n11335), .B1(n6183), .Y(n6594) );
  OAI22X1TS U6063 ( .A0(n10501), .A1(n10824), .B0(n10818), .B1(n10847), .Y(
        n6597) );
  AOI211X1TS U6060 ( .A0(n5798), .A1(n5314), .B0(n6591), .C0(n6592), .Y(n5404)
         );
  AOI22X1TS U6059 ( .A0(n10951), .A1(n6183), .B0(n10245), .B1(n6162), .Y(n6589) );
  AOI22X1TS U6057 ( .A0(n11343), .A1(n9993), .B0(n11669), .B1(n5617), .Y(n6590) );
  OAI211X1TS U6056 ( .A0(n10416), .A1(n10846), .B0(n6589), .C0(n6590), .Y(
        n6588) );
  OAI31X1TS U6054 ( .A0(n10716), .A1(n9432), .A2(n10985), .B0(n6586), .Y(n5787) );
  AOI22X1TS U6052 ( .A0(n10246), .A1(n6584), .B0(n11674), .B1(n6187), .Y(n6545) );
  AOI22X1TS U6051 ( .A0(n10145), .A1(n5807), .B0(n10555), .B1(n5783), .Y(n6546) );
  NOR3X1TS U6050 ( .A(n6583), .B(n10980), .C(n10044), .Y(n6186) );
  AOI211X1TS U6047 ( .A0(n9989), .A1(n6581), .B0(n6186), .C0(n6582), .Y(n6547)
         );
  NOR2X1TS U6046 ( .A(n12441), .B(n10185), .Y(n6549) );
  OAI211X1TS U6042 ( .A0(n10984), .A1(n10190), .B0(n6576), .C0(n6577), .Y(
        n5812) );
  OAI22X1TS U6040 ( .A0(n9312), .A1(n10521), .B0(n12494), .B1(n11672), .Y(
        n6550) );
  NOR2X1TS U6035 ( .A(n11684), .B(n10555), .Y(n5809) );
  AOI211X1TS U6032 ( .A0(n11670), .A1(n6011), .B0(n6570), .C0(n6571), .Y(n6568) );
  NOR2X1TS U6028 ( .A(n10189), .B(n11977), .Y(n5637) );
  AOI211X1TS U6024 ( .A0(n10558), .A1(n11397), .B0(n6561), .C0(n6562), .Y(
        n6559) );
  OAI211X1TS U6023 ( .A0(n6558), .A1(n12440), .B0(n6559), .C0(n6560), .Y(n6557) );
  AOI211X1TS U6022 ( .A0(n11696), .A1(n11377), .B0(n5618), .C0(n6557), .Y(
        n5403) );
  AOI22X1TS U6020 ( .A0(n11379), .A1(n9283), .B0(n11229), .B1(n6011), .Y(n6552) );
  NOR2X1TS U6010 ( .A(n11342), .B(n10953), .Y(n6189) );
  OAI22X1TS U5992 ( .A0(n12497), .A1(n10149), .B0(n11690), .B1(n9942), .Y(
        n6533) );
  NOR3X1TS U5991 ( .A(n6531), .B(n6532), .C(n6533), .Y(n5811) );
  INVX2TS U5983 ( .A(n5232), .Y(n5231) );
  NOR2X1TS U4636 ( .A(n12269), .B(n10917), .Y(n4392) );
  AOI22X1TS U4615 ( .A0(n11358), .A1(n11744), .B0(n12261), .B1(n11370), .Y(
        n4997) );
  OAI211X1TS U4614 ( .A0(n4392), .A1(n11262), .B0(n4996), .C0(n4997), .Y(n4995) );
  NOR2X1TS U4608 ( .A(n10109), .B(n10425), .Y(n4028) );
  AOI211X1TS U4587 ( .A0(n12259), .A1(n10451), .B0(n4990), .C0(n4991), .Y(
        n4989) );
  AOI211X1TS U4584 ( .A0(n12586), .A1(n10136), .B0(n4028), .C0(n4988), .Y(
        n3859) );
  AOI21X1TS U4576 ( .A0(n10140), .A1(n9666), .B0(n12443), .Y(n4622) );
  AOI22X1TS U4569 ( .A0(n11369), .A1(n12000), .B0(n11232), .B1(n11750), .Y(
        n4984) );
  OAI21X1TS U4568 ( .A0(n11340), .A1(n11363), .B0(n4984), .Y(n4983) );
  AOI211X1TS U4547 ( .A0(n11368), .A1(n3719), .B0(n4978), .C0(n4979), .Y(n4163) );
  NOR2X1TS U4517 ( .A(n3701), .B(n10767), .Y(n4031) );
  AOI211X1TS U4506 ( .A0(n11231), .A1(n12260), .B0(n3720), .C0(n4054), .Y(
        n4963) );
  OAI22X1TS U4503 ( .A0(n10398), .A1(n10394), .B0(n10481), .B1(n12009), .Y(
        n4958) );
  OAI22X1TS U4500 ( .A0(n4419), .A1(n10378), .B0(n3707), .B1(n11346), .Y(n4959) );
  OAI22X1TS U4497 ( .A0(n11351), .A1(n12010), .B0(n9138), .B1(n11345), .Y(
        n4957) );
  OAI211X1TS U4495 ( .A0(n9102), .A1(n12445), .B0(n4164), .C0(n4165), .Y(n4941) );
  NOR2X1TS U4494 ( .A(n11232), .B(n10450), .Y(n4064) );
  NOR2X1TS U4487 ( .A(n10405), .B(n12587), .Y(n4065) );
  OAI22X1TS U4484 ( .A0(n10377), .A1(n10399), .B0(n10139), .B1(n10839), .Y(
        n4949) );
  OAI22X1TS U4483 ( .A0(n10485), .A1(n11362), .B0(n10426), .B1(n12010), .Y(
        n4950) );
  NOR2X1TS U4482 ( .A(n10494), .B(n9906), .Y(n4588) );
  OAI22X1TS U5032 ( .A0(n12492), .A1(n10143), .B0(n12569), .B1(n12531), .Y(
        n5057) );
  OAI31X1TS U5024 ( .A0(n9788), .A1(n9196), .A2(n12538), .B0(n4560), .Y(n5058)
         );
  NOR2X1TS U5011 ( .A(n9922), .B(n10456), .Y(n4533) );
  AOI32X1TS U4993 ( .A0(n10860), .A1(n5114), .A2(n12531), .B0(n4492), .B1(
        n5114), .Y(n5113) );
  AOI211X1TS U4992 ( .A0(n9686), .A1(n10807), .B0(n4533), .C0(n5113), .Y(n4313) );
  AOI22X1TS U4981 ( .A0(n10147), .A1(n10808), .B0(n10133), .B1(n9098), .Y(
        n5107) );
  INVX2TS U4975 ( .A(n4849), .Y(n4301) );
  AOI22X1TS U4970 ( .A0(n10414), .A1(n12032), .B0(n10806), .B1(n10459), .Y(
        n5109) );
  OAI211X1TS U4966 ( .A0(n12533), .A1(n10143), .B0(n5109), .C0(n4870), .Y(
        n4318) );
  AOI211X1TS U4965 ( .A0(n10875), .A1(n10812), .B0(n4301), .C0(n4318), .Y(
        n5108) );
  NOR2X1TS U4960 ( .A(n9639), .B(n9651), .Y(n5076) );
  AOI211X1TS U4948 ( .A0(n10400), .A1(n11769), .B0(n4824), .C0(n5105), .Y(
        n5104) );
  OAI211X1TS U4946 ( .A0(n12207), .A1(n10776), .B0(n5104), .C0(n4547), .Y(
        n4317) );
  OAI22X1TS U4940 ( .A0(n9937), .A1(n10771), .B0(n10112), .B1(n12533), .Y(
        n5077) );
  NOR2X1TS U4936 ( .A(n10147), .B(n9687), .Y(n4573) );
  AOI22X1TS U4932 ( .A0(n10414), .A1(n4325), .B0(n10460), .B1(n4307), .Y(n5080) );
  AOI21X1TS U4930 ( .A0(n10112), .A1(n11773), .B0(n11715), .Y(n4576) );
  AOI211X1TS U4924 ( .A0(n10803), .A1(n4819), .B0(n4576), .C0(n5100), .Y(n5081) );
  NOR2X1TS U4911 ( .A(n11212), .B(n10414), .Y(n4319) );
  AOI21X1TS U4892 ( .A0(n12202), .A1(n10803), .B0(n5085), .Y(n4312) );
  NOR2X1TS U4881 ( .A(n11248), .B(n10807), .Y(n3962) );
  OAI22X1TS U4876 ( .A0(n10783), .A1(n11757), .B0(n12572), .B1(n11773), .Y(
        n5066) );
  AOI21X1TS U4874 ( .A0(n12571), .A1(n12530), .B0(n11763), .Y(n5068) );
  AOI22X1TS U4873 ( .A0(n10391), .A1(n4568), .B0(n10876), .B1(n4850), .Y(n5070) );
  NOR2X1TS U4868 ( .A(n11250), .B(n10395), .Y(n4320) );
  OAI22X1TS U4867 ( .A0(n4834), .A1(n12023), .B0(n4320), .B1(n10776), .Y(n5062) );
  NOR2X1TS U4866 ( .A(n11767), .B(n11702), .Y(n3967) );
  NOR2X1TS U4864 ( .A(n10115), .B(n12621), .Y(n3963) );
  AOI22X1TS U4184 ( .A0(n10882), .A1(n9917), .B0(n10370), .B1(n10160), .Y(
        n4793) );
  AOI22X1TS U4181 ( .A0(n11417), .A1(n4780), .B0(n11272), .B1(n4379), .Y(n4794) );
  AOI211X1TS U4177 ( .A0(n4013), .A1(n3516), .B0(n4791), .C0(n4792), .Y(n3606)
         );
  AOI22X1TS U4176 ( .A0(n10799), .A1(n4379), .B0(n10386), .B1(n4358), .Y(n4789) );
  OAI211X1TS U4173 ( .A0(n10499), .A1(n10921), .B0(n4789), .C0(n4790), .Y(
        n4788) );
  OAI31X1TS U4171 ( .A0(n10753), .A1(n9232), .A2(n10759), .B0(n4786), .Y(n4003) );
  AOI22X1TS U4169 ( .A0(n10386), .A1(n4784), .B0(n11785), .B1(n4383), .Y(n4745) );
  AOI22X1TS U4168 ( .A0(n10155), .A1(n4021), .B0(n10370), .B1(n3989), .Y(n4746) );
  NOR3X1TS U4167 ( .A(n4783), .B(n10764), .C(n10747), .Y(n4382) );
  AOI22X1TS U4166 ( .A0(n9180), .A1(n10126), .B0(n10434), .B1(n10881), .Y(
        n3510) );
  AOI211X1TS U4164 ( .A0(n9933), .A1(n4781), .B0(n4382), .C0(n4782), .Y(n4747)
         );
  NOR2X1TS U4163 ( .A(n12389), .B(n10123), .Y(n4749) );
  OAI211X1TS U4159 ( .A0(n10758), .A1(n10120), .B0(n4776), .C0(n4777), .Y(
        n3980) );
  AOI211X1TS U4155 ( .A0(n10385), .A1(n11809), .B0(n4774), .C0(n4775), .Y(
        n4766) );
  NOR2X1TS U4152 ( .A(n11797), .B(n10370), .Y(n3977) );
  INVX2TS U4151 ( .A(n3977), .Y(n4244) );
  NOR2X1TS U4147 ( .A(n10403), .B(n9665), .Y(n3823) );
  NOR2X1TS U4145 ( .A(n10119), .B(n12038), .Y(n3842) );
  AOI211X1TS U4141 ( .A0(n10374), .A1(n11220), .B0(n4761), .C0(n4762), .Y(
        n4759) );
  OAI211X1TS U4140 ( .A0(n4758), .A1(n12388), .B0(n4759), .C0(n4760), .Y(n4757) );
  AOI211X1TS U4139 ( .A0(n12072), .A1(n10784), .B0(n3823), .C0(n4757), .Y(
        n3605) );
  AOI22X1TS U4137 ( .A0(n10786), .A1(n9095), .B0(n10883), .B1(n4244), .Y(n4752) );
  NOR2X1TS U4127 ( .A(n11268), .B(n10801), .Y(n4386) );
  NOR2X1TS U4126 ( .A(n10130), .B(n10121), .Y(n3985) );
  OAI22X1TS U4120 ( .A0(n9122), .A1(n10788), .B0(n3846), .B1(n9919), .Y(n4741)
         );
  AOI22X1TS U4118 ( .A0(n10380), .A1(n10160), .B0(n10429), .B1(n9096), .Y(
        n4725) );
  OAI22X1TS U4112 ( .A0(n12388), .A1(n12548), .B0(n11709), .B1(n10152), .Y(
        n4728) );
  NOR3X1TS U4108 ( .A(n4731), .B(n4732), .C(n4733), .Y(n3979) );
  NOR4BX1TS U4103 ( .AN(n3606), .B(n4003), .C(n4230), .D(n4723), .Y(n3386) );
  INVX2TS U4100 ( .A(n3435), .Y(n3434) );
  OAI22X1TS U7446 ( .A0(n7681), .A1(n10661), .B0(n7850), .B1(n11867), .Y(n7840) );
  OAI211X1TS U7445 ( .A0(n7690), .A1(n9552), .B0(n7848), .C0(n7849), .Y(n7841)
         );
  OAI211X1TS U7443 ( .A0(n11611), .A1(n11920), .B0(n7844), .C0(n7845), .Y(
        n7842) );
  OAI22X1TS U7438 ( .A0(n7833), .A1(n10343), .B0(n7834), .B1(n11922), .Y(n7832) );
  OAI211X1TS U7428 ( .A0(n11107), .A1(n11904), .B0(n7813), .C0(n7814), .Y(
        n7812) );
  AOI211X1TS U7427 ( .A0(n10282), .A1(n7810), .B0(n7811), .C0(n7812), .Y(n7809) );
  INVX2TS U7425 ( .A(n9216), .Y(n6943) );
  AOI22X1TS U6955 ( .A0(n6943), .A1(n1605), .B0(n1607), .B1(n9216), .Y(n6939)
         );
  INVX2TS U7027 ( .A(n1298), .Y(n1297) );
  AOI22X1TS U8312 ( .A0(n12627), .A1(n8529), .B0(n10090), .B1(n7979), .Y(n8527) );
  AOI22X1TS U8310 ( .A0(n10102), .A1(n11194), .B0(n12596), .B1(n8529), .Y(
        n8528) );
  OAI211X1TS U8309 ( .A0(n10697), .A1(n12163), .B0(n8527), .C0(n8528), .Y(
        n8526) );
  AOI211X1TS U8308 ( .A0(n11493), .A1(n8219), .B0(n8397), .C0(n8526), .Y(n8524) );
  AOI22X1TS U8301 ( .A0(n11579), .A1(n10638), .B0(n11092), .B1(n7610), .Y(
        n8513) );
  AOI211X1TS U8282 ( .A0(n11581), .A1(n9531), .B0(n8248), .C0(n8515), .Y(n8514) );
  OAI211X1TS U8281 ( .A0(n10094), .A1(n11164), .B0(n8513), .C0(n8514), .Y(
        n8512) );
  OAI22X1TS U8277 ( .A0(n8413), .A1(n11892), .B0(n8179), .B1(n10050), .Y(n8480) );
  OAI31X1TS U8264 ( .A0(n10333), .A1(n11503), .A2(n7451), .B0(n12481), .Y(
        n8504) );
  OAI211X1TS U8263 ( .A0(n8503), .A1(n10097), .B0(n7469), .C0(n8504), .Y(n8481) );
  AOI211X1TS U8237 ( .A0(n11492), .A1(n12635), .B0(n8227), .C0(n8489), .Y(
        n8483) );
  OAI22X1TS U8233 ( .A0(n11892), .A1(n11952), .B0(n12171), .B1(n12128), .Y(
        n8487) );
  AOI211X1TS U8232 ( .A0(n11944), .A1(n9511), .B0(n8486), .C0(n8487), .Y(n8485) );
  NOR4BX1TS U8230 ( .AN(n7957), .B(n8480), .C(n8481), .D(n8482), .Y(n6980) );
  OAI22X1TS U8034 ( .A0(n9128), .A1(n9213), .B0(n7028), .B1(n6980), .Y(n1279)
         );
  INVX2TS U8033 ( .A(n1279), .Y(n1276) );
  AOI22X1TS U1142 ( .A0(n1297), .A1(n12661), .B0(n1279), .B1(n1298), .Y(n1290)
         );
  AOI221X1TS U7970 ( .A0(n11580), .A1(n12643), .B0(n10701), .B1(n12471), .C0(
        n8362), .Y(n7627) );
  OAI32X1TS U7958 ( .A0(n8353), .A1(n11946), .A2(n11581), .B0(n12597), .B1(
        n8353), .Y(n8352) );
  OAI211X1TS U7956 ( .A0(n11198), .A1(n11575), .B0(n8352), .C0(n7463), .Y(
        n7576) );
  OAI22X1TS U1137 ( .A0(n1288), .A1(n12764), .B0(n12692), .B1(n1289), .Y(N97)
         );
  AOI22X1TS U7548 ( .A0(n10702), .A1(n7451), .B0(n10692), .B1(n9486), .Y(n7966) );
  AOI211X1TS U7546 ( .A0(n10310), .A1(n9822), .B0(n7961), .C0(n7962), .Y(n7958) );
  NOR4BX1TS U7543 ( .AN(n7954), .B(n7955), .C(n7444), .D(n7956), .Y(n6923) );
  INVX2TS U7371 ( .A(n6923), .Y(n1645) );
  AOI211X1TS U7369 ( .A0(n11138), .A1(n11927), .B0(n7740), .C0(n7741), .Y(
        n7735) );
  OAI22X1TS U7368 ( .A0(n10656), .A1(n11867), .B0(n9846), .B1(n10718), .Y(
        n7738) );
  AOI221X1TS U7367 ( .A0(n12633), .A1(n11155), .B0(n12184), .B1(n11862), .C0(
        n7738), .Y(n7736) );
  OAI211X1TS U7366 ( .A0(n10724), .A1(n10029), .B0(n7735), .C0(n7736), .Y(
        n7706) );
  AOI32X1TS U7353 ( .A0(n7714), .A1(n11922), .A2(n9492), .B0(n10713), .B1(
        n7714), .Y(n7713) );
  AOI211X1TS U7352 ( .A0(n11915), .A1(n7712), .B0(n7697), .C0(n7713), .Y(n7709) );
  OAI31X1TS U7351 ( .A0(n12364), .A1(n11854), .A2(n10069), .B0(n12351), .Y(
        n7710) );
  INVX2TS U7346 ( .A(n6986), .Y(n6985) );
  AOI22X1TS U7511 ( .A0(n10270), .A1(n7797), .B0(n11050), .B1(n7074), .Y(n7918) );
  AOI22X1TS U7510 ( .A0(n10674), .A1(n9801), .B0(n10591), .B1(n7920), .Y(n7919) );
  OAI211X1TS U7509 ( .A0(n10618), .A1(n10010), .B0(n7918), .C0(n7919), .Y(
        n7917) );
  AOI211X1TS U7508 ( .A0(n11886), .A1(n7171), .B0(n7441), .C0(n7917), .Y(n7909) );
  OAI211X1TS U7502 ( .A0(n7432), .A1(n11796), .B0(n7909), .C0(n7910), .Y(n7908) );
  NOR2X1TS U6714 ( .A(n12243), .B(n10870), .Y(n6235) );
  AOI22X1TS U6693 ( .A0(n11293), .A1(n11704), .B0(n12250), .B1(n11283), .Y(
        n6854) );
  OAI211X1TS U6692 ( .A0(n6235), .A1(n11367), .B0(n6853), .C0(n6854), .Y(n6852) );
  NOR2X1TS U6686 ( .A(n10221), .B(n10512), .Y(n5884) );
  AOI211X1TS U6665 ( .A0(n12247), .A1(n10465), .B0(n6847), .C0(n6848), .Y(
        n6846) );
  AOI211X1TS U6662 ( .A0(n12590), .A1(n10170), .B0(n5884), .C0(n6845), .Y(
        n5714) );
  AOI21X1TS U6654 ( .A0(n10166), .A1(n9706), .B0(n12399), .Y(n6494) );
  AOI22X1TS U6647 ( .A0(n11282), .A1(n12048), .B0(n11415), .B1(n11698), .Y(
        n6841) );
  OAI21X1TS U6646 ( .A0(n11312), .A1(n11288), .B0(n6841), .Y(n6840) );
  OAI22X1TS U6631 ( .A0(n10221), .A1(n10537), .B0(n10448), .B1(n10918), .Y(
        n6835) );
  AOI211X1TS U6625 ( .A0(n11281), .A1(n5540), .B0(n6835), .C0(n6836), .Y(n6117) );
  NOR2X1TS U6595 ( .A(n12273), .B(n11013), .Y(n5887) );
  AOI211X1TS U6584 ( .A0(n11413), .A1(n12248), .B0(n5541), .C0(n5910), .Y(
        n6820) );
  OAI22X1TS U6581 ( .A0(n10537), .A1(n10542), .B0(n10453), .B1(n12041), .Y(
        n6815) );
  OAI22X1TS U6578 ( .A0(n6262), .A1(n10573), .B0(n5528), .B1(n11307), .Y(n6816) );
  OAI22X1TS U6575 ( .A0(n11300), .A1(n12042), .B0(n9349), .B1(n11306), .Y(
        n6814) );
  NOR2X1TS U6572 ( .A(n11415), .B(n10466), .Y(n5920) );
  NOR2X1TS U6565 ( .A(n10586), .B(n5931), .Y(n5921) );
  OAI22X1TS U6562 ( .A0(n10572), .A1(n10536), .B0(n10165), .B1(n10931), .Y(
        n6806) );
  OAI22X1TS U6561 ( .A0(n10448), .A1(n11287), .B0(n10511), .B1(n12042), .Y(
        n6807) );
  NOR2X1TS U6560 ( .A(n10440), .B(n9962), .Y(n6460) );
  AOI22X1TS U5103 ( .A0(n9268), .A1(n5182), .B0(n9210), .B1(n5150), .Y(n5181)
         );
  AOI22X1TS U6991 ( .A0(n9456), .A1(n6976), .B0(n9224), .B1(n12678), .Y(n6975)
         );
  AOI22X1TS U5153 ( .A0(n9267), .A1(n5132), .B0(n9203), .B1(n5150), .Y(n5236)
         );
  NOR2X1TS U4831 ( .A(n12246), .B(n10899), .Y(n4432) );
  AOI22X1TS U4810 ( .A0(n11308), .A1(n11726), .B0(n12239), .B1(n11321), .Y(
        n5055) );
  OAI211X1TS U4809 ( .A0(n4432), .A1(n11255), .B0(n5054), .C0(n5055), .Y(n5053) );
  NOR2X1TS U4803 ( .A(n10117), .B(n10418), .Y(n4084) );
  AOI211X1TS U4782 ( .A0(n12237), .A1(n10443), .B0(n5048), .C0(n5049), .Y(
        n5047) );
  AOI211X1TS U4779 ( .A0(n12578), .A1(n10127), .B0(n4084), .C0(n5046), .Y(
        n3884) );
  AOI21X1TS U4771 ( .A0(n10132), .A1(n9662), .B0(n12427), .Y(n4694) );
  AOI22X1TS U4764 ( .A0(n11322), .A1(n11987), .B0(n11225), .B1(n11731), .Y(
        n5042) );
  OAI21X1TS U4763 ( .A0(n11291), .A1(n11315), .B0(n5042), .Y(n5041) );
  OAI22X1TS U4748 ( .A0(n10117), .A1(n10389), .B0(n10467), .B1(n10821), .Y(
        n5036) );
  AOI211X1TS U4742 ( .A0(n11320), .A1(n3785), .B0(n5036), .C0(n5037), .Y(n4207) );
  NOR2X1TS U4712 ( .A(n12214), .B(n10780), .Y(n4087) );
  AOI211X1TS U4701 ( .A0(n11225), .A1(n12239), .B0(n3786), .C0(n4110), .Y(
        n5021) );
  OAI22X1TS U4698 ( .A0(n10388), .A1(n10383), .B0(n10464), .B1(n11994), .Y(
        n5016) );
  OAI22X1TS U4695 ( .A0(n4459), .A1(n10373), .B0(n3773), .B1(n11298), .Y(n5017) );
  OAI22X1TS U4692 ( .A0(n11303), .A1(n11995), .B0(n9150), .B1(n11297), .Y(
        n5015) );
  NOR2X1TS U4689 ( .A(n11226), .B(n10442), .Y(n4120) );
  NOR2X1TS U4682 ( .A(n10408), .B(n12578), .Y(n4121) );
  OAI22X1TS U4679 ( .A0(n10373), .A1(n10387), .B0(n10132), .B1(n10811), .Y(
        n5007) );
  OAI22X1TS U4678 ( .A0(n10467), .A1(n11314), .B0(n10420), .B1(n11995), .Y(
        n5008) );
  NOR2X1TS U4677 ( .A(n10476), .B(n9910), .Y(n4660) );
  INVX2TS U3272 ( .A(n9081), .Y(n3353) );
  AOI22X1TS U3223 ( .A0(n3353), .A1(n3386), .B0(n9195), .B1(n9080), .Y(n3385)
         );
  NOR2X1TS U3768 ( .A(n9913), .B(n10108), .Y(n3621) );
  NOR2X1TS U3767 ( .A(n10764), .B(n9930), .Y(n4248) );
  AOI211X1TS U3766 ( .A0(n10385), .A1(n9918), .B0(n3621), .C0(n4248), .Y(n4353) );
  AOI31X1TS U3765 ( .A0(n12388), .A1(n9664), .A2(n11388), .B0(n12549), .Y(
        n4355) );
  AOI211X1TS U3762 ( .A0(n10933), .A1(n11219), .B0(n4355), .C0(n4356), .Y(
        n4354) );
  OAI22X1TS U3462 ( .A0(n3837), .A1(n4273), .B0(n12037), .B1(n10795), .Y(n3824) );
  OAI22X1TS U3461 ( .A0(n3613), .A1(n3841), .B0(n9914), .B1(n11387), .Y(n3825)
         );
  AOI32X1TS U3340 ( .A0(n3515), .A1(n4256), .A2(n3517), .B0(n10921), .B1(n3515), .Y(n3505) );
  OAI211X1TS U3338 ( .A0(n3507), .A1(n12275), .B0(n3509), .C0(n3510), .Y(n3506) );
  AOI211X1TS U3337 ( .A0(n10934), .A1(n9095), .B0(n3505), .C0(n3506), .Y(n3480) );
  OAI22X1TS U3336 ( .A0(n12548), .A1(n11803), .B0(n12283), .B1(n10152), .Y(
        n3483) );
  OAI22X1TS U3335 ( .A0(n10504), .A1(n12064), .B0(n10938), .B1(n9920), .Y(
        n3484) );
  NOR2X1TS U3692 ( .A(n11388), .B(n10124), .Y(n3494) );
  AOI221X1TS U3334 ( .A0(n11809), .A1(n10159), .B0(n12074), .B1(n10156), .C0(
        n3494), .Y(n3488) );
  OAI22X1TS U3784 ( .A0(n10943), .A1(n11388), .B0(n12276), .B1(n10124), .Y(
        n4374) );
  INVX2TS U3781 ( .A(n9121), .Y(n3990) );
  AOI22X1TS U3271 ( .A0(n3353), .A1(n3340), .B0(n1555), .B1(n9081), .Y(n3439)
         );
  INVX2TS U8422 ( .A(n6952), .Y(n6951) );
  OAI22X1TS U7814 ( .A0(n8221), .A1(n12733), .B0(n12683), .B1(n8222), .Y(N100)
         );
  AOI22X1TS U4071 ( .A0(n10409), .A1(n3887), .B0(n11727), .B1(n4698), .Y(n4668) );
  OAI22X1TS U4067 ( .A0(n4660), .A1(n11302), .B0(n9655), .B1(n12397), .Y(n4206) );
  OAI211X1TS U4045 ( .A0(n3805), .A1(n9162), .B0(n4674), .C0(n4675), .Y(n4673)
         );
  NOR4BX1TS U4044 ( .AN(n4671), .B(n3778), .C(n4672), .D(n4673), .Y(n4670) );
  AOI22X1TS U4034 ( .A0(n12580), .A1(n10827), .B0(n11278), .B1(n9114), .Y(
        n3890) );
  OAI22X1TS U4033 ( .A0(n11303), .A1(n11256), .B0(n9147), .B1(n12430), .Y(
        n4657) );
  NOR4BX1TS U4030 ( .AN(n3890), .B(n4657), .C(n4658), .D(n4659), .Y(n4652) );
  AOI221X1TS U4027 ( .A0(n10443), .A1(n9186), .B0(n11733), .B1(n12053), .C0(
        n4655), .Y(n4654) );
  NOR4BX1TS U4025 ( .AN(n3741), .B(n3779), .C(n4101), .D(n4651), .Y(n1584) );
  AOI22X1TS U3996 ( .A0(n10404), .A1(n3862), .B0(n11745), .B1(n4626), .Y(n4596) );
  OAI22X1TS U3992 ( .A0(n4588), .A1(n11350), .B0(n9659), .B1(n12404), .Y(n4162) );
  OAI211X1TS U3970 ( .A0(n3739), .A1(n9154), .B0(n4602), .C0(n4603), .Y(n4601)
         );
  NOR4BX1TS U3969 ( .AN(n4599), .B(n3712), .C(n4600), .D(n4601), .Y(n4598) );
  AOI22X1TS U3959 ( .A0(n12585), .A1(n10855), .B0(n11326), .B1(n9106), .Y(
        n3865) );
  NOR4BX1TS U3955 ( .AN(n3865), .B(n4585), .C(n4586), .D(n4587), .Y(n4580) );
  NOR4BX1TS U3950 ( .AN(n3675), .B(n3713), .C(n4045), .D(n4579), .Y(n1626) );
  NOR2X1TS U3867 ( .A(n10805), .B(n11284), .Y(n3891) );
  OAI22X1TS U3865 ( .A0(n3891), .A1(n12398), .B0(n3589), .B1(n10418), .Y(n4455) );
  AOI22X1TS U3861 ( .A0(n12507), .A1(n9909), .B0(n10780), .B1(n9642), .Y(n4460) );
  OAI22X1TS U3858 ( .A0(n10371), .A1(n9663), .B0(n10437), .B1(n11291), .Y(
        n4447) );
  OAI22X1TS U3857 ( .A0(n3788), .A1(n10382), .B0(n11315), .B1(n12430), .Y(
        n4448) );
  AOI211X1TS U3855 ( .A0(n10477), .A1(n11286), .B0(n4452), .C0(n4453), .Y(
        n4451) );
  OAI211X1TS U3854 ( .A0(n10131), .A1(n10113), .B0(n4450), .C0(n4451), .Y(
        n4449) );
  OAI22X1TS U3852 ( .A0(n11398), .A1(n12429), .B0(n9663), .B1(n11236), .Y(
        n4440) );
  OAI22X1TS U3851 ( .A0(n11256), .A1(n10894), .B0(n10373), .B1(n10418), .Y(
        n4441) );
  OAI21X1TS U3850 ( .A0(n12238), .A1(n10772), .B0(n10779), .Y(n4445) );
  OAI211X1TS U3848 ( .A0(n12428), .A1(n10821), .B0(n4445), .C0(n3764), .Y(
        n4442) );
  AOI31X1TS U3844 ( .A0(n9111), .A1(n11398), .A2(n10893), .B0(n11996), .Y(
        n4428) );
  AOI21X1TS U3843 ( .A0(n9186), .A1(n9144), .B0(n11393), .Y(n4224) );
  OAI22X1TS U3842 ( .A0(n9110), .A1(n9672), .B0(n4224), .B1(n11304), .Y(n4430)
         );
  AOI22X1TS U3841 ( .A0(n4203), .A1(n4119), .B0(n11308), .B1(n9165), .Y(n4433)
         );
  OAI211X1TS U3835 ( .A0(n4432), .A1(n3802), .B0(n4433), .C0(n4434), .Y(n4431)
         );
  NOR2X1TS U3900 ( .A(n9118), .B(n10397), .Y(n3916) );
  AOI22X1TS U3897 ( .A0(n9175), .A1(n4513), .B0(n10877), .B1(n4306), .Y(n4510)
         );
  OAI211X1TS U3895 ( .A0(n4509), .A1(n10860), .B0(n4510), .C0(n4511), .Y(n4508) );
  AOI211X1TS U3894 ( .A0(n10807), .A1(n9680), .B0(n4507), .C0(n4508), .Y(n4505) );
  OAI211X1TS U3893 ( .A0(n3916), .A1(n12540), .B0(n4504), .C0(n4505), .Y(n4287) );
  AOI22X1TS U3891 ( .A0(n10814), .A1(n4502), .B0(n11375), .B1(n10133), .Y(
        n4494) );
  OAI22X1TS U3889 ( .A0(n12490), .A1(n10792), .B0(n10871), .B1(n10112), .Y(
        n4500) );
  NOR2X1TS U3947 ( .A(n10797), .B(n10415), .Y(n3910) );
  OAI22X1TS U3879 ( .A0(n11761), .A1(n9676), .B0(n11773), .B1(n12023), .Y(
        n4477) );
  AOI22X1TS U3878 ( .A0(n9176), .A1(n3668), .B0(n12619), .B1(n10134), .Y(n4479) );
  OAI211X1TS U3876 ( .A0(n10144), .A1(n10776), .B0(n4479), .C0(n3661), .Y(
        n4478) );
  AOI211X1TS U3875 ( .A0(n10148), .A1(n11213), .B0(n4477), .C0(n4478), .Y(
        n4469) );
  OAI22X1TS U3872 ( .A0(n4474), .A1(n11763), .B0(n9937), .B1(n12493), .Y(n4473) );
  OAI31X1TS U3870 ( .A0(n9118), .A1(n11702), .A2(n9099), .B0(n12030), .Y(n4471) );
  NOR2X1TS U3716 ( .A(n9904), .B(n10130), .Y(n3618) );
  OAI211X1TS U3711 ( .A0(n4276), .A1(n10755), .B0(n4277), .C0(n4278), .Y(n4275) );
  AOI211X1TS U3710 ( .A0(n10379), .A1(n10385), .B0(n4274), .C0(n4275), .Y(
        n4271) );
  OAI211X1TS U3709 ( .A0(n3618), .A1(n12065), .B0(n4270), .C0(n4271), .Y(n4004) );
  OAI22X1TS U3708 ( .A0(n10499), .A1(n3511), .B0(n12389), .B1(n10765), .Y(
        n4264) );
  NOR2X1TS U3794 ( .A(n10370), .B(n11785), .Y(n3612) );
  OAI22X1TS U3707 ( .A0(n3612), .A1(n10498), .B0(n12282), .B1(n11387), .Y(
        n4265) );
  NOR2X1TS U3706 ( .A(n4272), .B(n10123), .Y(n3816) );
  OAI211X1TS U3703 ( .A0(n10943), .A1(n10164), .B0(n4267), .C0(n4268), .Y(
        n4266) );
  OAI22X1TS U3701 ( .A0(n12390), .A1(n10787), .B0(n12277), .B1(n10793), .Y(
        n4249) );
  AOI22X1TS U3698 ( .A0(n10374), .A1(n10122), .B0(n10785), .B1(n10125), .Y(
        n4254) );
  OAI22X1TS U3695 ( .A0(n4247), .A1(n10503), .B0(n9121), .B1(n11708), .Y(n4234) );
  AOI211X1TS U3687 ( .A0(n11267), .A1(n9096), .B0(n4234), .C0(n4235), .Y(n4232) );
  NOR3X1TS U3684 ( .A(n4004), .B(n4230), .C(n4231), .Y(n3372) );
  AOI22X1TS U3253 ( .A0(n3420), .A1(n3421), .B0(n3422), .B1(n12657), .Y(n3419)
         );
  INVX2TS U3265 ( .A(n3408), .Y(n3407) );
  AOI22X1TS U3264 ( .A0(n3433), .A1(n3434), .B0(n3435), .B1(n1583), .Y(n3432)
         );
  AOI22X1TS U7000 ( .A0(n6984), .A1(n6985), .B0(n6986), .B1(n1567), .Y(n6983)
         );
  AOI22X1TS U7055 ( .A0(n6943), .A1(n6985), .B0(n6986), .B1(n9217), .Y(n7031)
         );
  NOR2X1TS U3831 ( .A(n10833), .B(n11333), .Y(n3866) );
  OAI22X1TS U3829 ( .A0(n3866), .A1(n12404), .B0(n3550), .B1(n10424), .Y(n4415) );
  AOI22X1TS U3827 ( .A0(n12260), .A1(n12058), .B0(n11328), .B1(n10768), .Y(
        n4423) );
  AOI22X1TS U3825 ( .A0(n12523), .A1(n9905), .B0(n10767), .B1(n9646), .Y(n4420) );
  OAI211X1TS U3824 ( .A0(n4419), .A1(n11261), .B0(n4420), .C0(n4421), .Y(n4418) );
  OAI22X1TS U3822 ( .A0(n10376), .A1(n9667), .B0(n10447), .B1(n11339), .Y(
        n4407) );
  OAI22X1TS U3821 ( .A0(n3722), .A1(n10393), .B0(n11364), .B1(n12443), .Y(
        n4408) );
  AOI211X1TS U3819 ( .A0(n10493), .A1(n11334), .B0(n4412), .C0(n4413), .Y(
        n4411) );
  OAI211X1TS U3818 ( .A0(n10140), .A1(n10105), .B0(n4410), .C0(n4411), .Y(
        n4409) );
  OAI22X1TS U3816 ( .A0(n11410), .A1(n12446), .B0(n9666), .B1(n11243), .Y(
        n4400) );
  OAI22X1TS U3815 ( .A0(n11260), .A1(n10911), .B0(n10378), .B1(n10426), .Y(
        n4401) );
  OAI21X1TS U3814 ( .A0(n12259), .A1(n10760), .B0(n10766), .Y(n4405) );
  OAI211X1TS U3812 ( .A0(n12444), .A1(n10850), .B0(n4405), .C0(n3698), .Y(
        n4402) );
  AOI31X1TS U3808 ( .A0(n9103), .A1(n11410), .A2(n10910), .B0(n3693), .Y(n4388) );
  AOI21X1TS U3807 ( .A0(n9183), .A1(n9132), .B0(n11405), .Y(n4180) );
  OAI22X1TS U3806 ( .A0(n9102), .A1(n9669), .B0(n4180), .B1(n11352), .Y(n4390)
         );
  AOI22X1TS U3805 ( .A0(n12270), .A1(n10854), .B0(n11356), .B1(n9157), .Y(
        n4393) );
  OAI211X1TS U3799 ( .A0(n4392), .A1(n3736), .B0(n4393), .C0(n4394), .Y(n4391)
         );
  AOI22X1TS U3795 ( .A0(n9904), .A1(n10156), .B0(n11417), .B1(n10430), .Y(
        n4360) );
  AOI211X1TS U3787 ( .A0(n3500), .A1(n4383), .B0(n4384), .C0(n4385), .Y(n4380)
         );
  AOI211X1TS U3775 ( .A0(n11799), .A1(n11272), .B0(n4371), .C0(n4372), .Y(
        n4368) );
  AOI22X1TS U3770 ( .A0(n10155), .A1(n4358), .B0(n11811), .B1(n3989), .Y(n4342) );
  OAI22X1TS U3757 ( .A0(n3837), .A1(n10403), .B0(n10151), .B1(n10795), .Y(
        n3608) );
  NOR3X1TS U3751 ( .A(n4339), .B(n3810), .C(n4340), .Y(n1546) );
  INVX2TS U5147 ( .A(n5205), .Y(n5204) );
  AOI22X1TS U5146 ( .A0(n5230), .A1(n5231), .B0(n5232), .B1(n1569), .Y(n5229)
         );
  NOR2X1TS U2929 ( .A(n2430), .B(n9282), .Y(n2864) );
  NOR2X1TS U2965 ( .A(n10322), .B(n10032), .Y(n3259) );
  AOI22X1TS U1794 ( .A0(n9971), .A1(n10199), .B0(n10248), .B1(n11870), .Y(
        n2441) );
  NOR2X1TS U2127 ( .A(n12367), .B(n10635), .Y(n2815) );
  INVX2TS U2094 ( .A(n2815), .Y(n2126) );
  NOR2X1TS U2947 ( .A(n9119), .B(n10028), .Y(n2723) );
  INVX2TS U2946 ( .A(n2723), .Y(n3250) );
  NOR2X1TS U1793 ( .A(n9980), .B(n10574), .Y(n1905) );
  NOR2X1TS U1792 ( .A(n11601), .B(n11471), .Y(n2259) );
  AOI211X1TS U1791 ( .A0(n10240), .A1(n2126), .B0(n1905), .C0(n2259), .Y(n2442) );
  NOR2X1TS U2101 ( .A(n11607), .B(n10997), .Y(n2455) );
  NOR2X1TS U2918 ( .A(n10700), .B(n2274), .Y(n3241) );
  NOR2X1TS U2021 ( .A(n9741), .B(n11567), .Y(n2239) );
  AOI22X1TS U2018 ( .A0(n10636), .A1(n11095), .B0(n12303), .B1(n10986), .Y(
        n2727) );
  OAI21X1TS U2017 ( .A0(n10200), .A1(n11131), .B0(n11115), .Y(n2728) );
  NOR2X1TS U2081 ( .A(n10219), .B(n11126), .Y(n2730) );
  NOR2X1TS U2016 ( .A(n9724), .B(n10296), .Y(n1763) );
  AOI211X1TS U1790 ( .A0(n10986), .A1(n10259), .B0(n2455), .C0(n2456), .Y(
        n2443) );
  NOR2X1TS U2857 ( .A(n10653), .B(n11882), .Y(n1917) );
  NOR2X1TS U2856 ( .A(n12467), .B(n10216), .Y(n2289) );
  AOI211X1TS U2855 ( .A0(n12303), .A1(n12604), .B0(n1917), .C0(n2289), .Y(
        n3234) );
  NOR2X1TS U2853 ( .A(n11601), .B(n11613), .Y(n2854) );
  NOR2X1TS U2895 ( .A(n10561), .B(n11924), .Y(n2725) );
  AOI211X1TS U2848 ( .A0(n10200), .A1(n12605), .B0(n2854), .C0(n3236), .Y(
        n3235) );
  AOI22X1TS U2832 ( .A0(n9627), .A1(n11084), .B0(n9972), .B1(n12301), .Y(n3220) );
  AOI22X1TS U2830 ( .A0(n11117), .A1(n12366), .B0(n10987), .B1(n9756), .Y(
        n3221) );
  NOR2X1TS U2829 ( .A(n11089), .B(n12303), .Y(n2279) );
  NOR2X1TS U2884 ( .A(n12130), .B(n11495), .Y(n2431) );
  NOR2X1TS U2827 ( .A(n2431), .B(n10998), .Y(n1929) );
  NOR2X1TS U2825 ( .A(n10199), .B(n11085), .Y(n2819) );
  OAI22X1TS U2824 ( .A0(n3225), .A1(n12087), .B0(n2819), .B1(n11614), .Y(n3224) );
  AOI211X1TS U2823 ( .A0(n11840), .A1(n3223), .B0(n1929), .C0(n3224), .Y(n3222) );
  AOI21X1TS U2007 ( .A0(n2723), .A1(n10323), .B0(n9948), .Y(n2449) );
  NOR2X1TS U2842 ( .A(n10565), .B(n11088), .Y(n2423) );
  OAI22X1TS U2129 ( .A0(n2272), .A1(n11607), .B0(n10992), .B1(n11601), .Y(
        n2102) );
  AOI22X1TS U1607 ( .A0(n11094), .A1(n2119), .B0(n11925), .B1(n2120), .Y(n2118) );
  NOR2X1TS U2968 ( .A(n11464), .B(n11127), .Y(n2798) );
  OAI211X1TS U2934 ( .A0(n12469), .A1(n11606), .B0(n2292), .C0(n2863), .Y(
        n3254) );
  NOR2X1TS U2920 ( .A(n11606), .B(n11120), .Y(n2268) );
  NOR2X1TS U2914 ( .A(n10992), .B(n10251), .Y(n2841) );
  AOI211X1TS U2913 ( .A0(n9947), .A1(n11084), .B0(n2268), .C0(n2841), .Y(n3257) );
  NOR2X1TS U2803 ( .A(n11613), .B(n10999), .Y(n2830) );
  NOR2X1TS U2873 ( .A(n12131), .B(n11930), .Y(n1931) );
  OAI22X1TS U2001 ( .A0(n12466), .A1(n12460), .B0(n10992), .B1(n12347), .Y(
        n2713) );
  AOI22X1TS U1998 ( .A0(n10579), .A1(n9058), .B0(n11871), .B1(n2719), .Y(n2717) );
  NOR2X1TS U2146 ( .A(n11875), .B(n10569), .Y(n2109) );
  NOR2X1TS U1694 ( .A(n11122), .B(n11883), .Y(n2114) );
  NOR2X1TS U1679 ( .A(n11573), .B(n9079), .Y(n2115) );
  AOI211X1TS U1605 ( .A0(n11094), .A1(n9757), .B0(n2114), .C0(n2115), .Y(n2111) );
  AOI32X1TS U1603 ( .A0(n10659), .A1(n2111), .A2(n1754), .B0(n12467), .B1(
        n2111), .Y(n2110) );
  AOI211X1TS U1602 ( .A0(n11090), .A1(n9627), .B0(n2109), .C0(n2110), .Y(n2108) );
  NOR2X1TS U2732 ( .A(n2386), .B(n9362), .Y(n2940) );
  NOR2X1TS U2768 ( .A(n10330), .B(n10064), .Y(n3199) );
  AOI22X1TS U1767 ( .A0(n9983), .A1(n10204), .B0(n10272), .B1(n11893), .Y(
        n2397) );
  NOR2X1TS U2202 ( .A(n12374), .B(n10645), .Y(n2891) );
  INVX2TS U2169 ( .A(n2891), .Y(n2100) );
  NOR2X1TS U2750 ( .A(n9123), .B(n10060), .Y(n2690) );
  INVX2TS U2749 ( .A(n2690), .Y(n3190) );
  NOR2X1TS U1766 ( .A(n9992), .B(n10547), .Y(n1842) );
  NOR2X1TS U1765 ( .A(n11620), .B(n11483), .Y(n2326) );
  AOI211X1TS U1764 ( .A0(n10264), .A1(n2100), .B0(n1842), .C0(n2326), .Y(n2398) );
  NOR2X1TS U2176 ( .A(n11624), .B(n10982), .Y(n2411) );
  NOR2X1TS U2721 ( .A(n10726), .B(n2341), .Y(n3181) );
  NOR2X1TS U1979 ( .A(n9745), .B(n2319), .Y(n2306) );
  AOI22X1TS U1976 ( .A0(n10644), .A1(n1845), .B0(n12297), .B1(n10973), .Y(
        n2694) );
  OAI21X1TS U1975 ( .A0(n10204), .A1(n11154), .B0(n11135), .Y(n2695) );
  NOR2X1TS U2156 ( .A(n10211), .B(n11147), .Y(n2697) );
  NOR2X1TS U1974 ( .A(n9728), .B(n10300), .Y(n1725) );
  AOI211X1TS U1763 ( .A0(n10971), .A1(n10283), .B0(n2411), .C0(n2412), .Y(
        n2399) );
  NOR2X1TS U2660 ( .A(n10667), .B(n11906), .Y(n1854) );
  NOR2X1TS U2659 ( .A(n12485), .B(n10207), .Y(n2356) );
  AOI211X1TS U2658 ( .A0(n12297), .A1(n12600), .B0(n1854), .C0(n2356), .Y(
        n3174) );
  NOR2X1TS U2656 ( .A(n11620), .B(n11630), .Y(n2930) );
  NOR2X1TS U2698 ( .A(n10533), .B(n11937), .Y(n2692) );
  AOI211X1TS U2651 ( .A0(n10204), .A1(n12601), .B0(n2930), .C0(n3176), .Y(
        n3175) );
  AOI22X1TS U2635 ( .A0(n9632), .A1(n11099), .B0(n9983), .B1(n12295), .Y(n3160) );
  NOR2X1TS U2632 ( .A(n11106), .B(n12297), .Y(n2346) );
  NOR2X1TS U2687 ( .A(n12147), .B(n11488), .Y(n2387) );
  NOR2X1TS U2630 ( .A(n2387), .B(n1880), .Y(n1866) );
  NOR2X1TS U2629 ( .A(n10528), .B(n10553), .Y(n3165) );
  NOR2X1TS U2628 ( .A(n10203), .B(n11100), .Y(n2895) );
  OAI22X1TS U2627 ( .A0(n3165), .A1(n12079), .B0(n2895), .B1(n11632), .Y(n3164) );
  AOI21X1TS U1965 ( .A0(n2690), .A1(n10331), .B0(n9944), .Y(n2405) );
  NOR2X1TS U2645 ( .A(n10539), .B(n11104), .Y(n2379) );
  OAI22X1TS U2204 ( .A0(n2339), .A1(n11625), .B0(n10977), .B1(n11619), .Y(
        n2076) );
  NOR2X1TS U2771 ( .A(n11477), .B(n11148), .Y(n2874) );
  OAI211X1TS U2737 ( .A0(n12483), .A1(n11624), .B0(n2359), .C0(n2939), .Y(
        n3194) );
  NOR2X1TS U2723 ( .A(n11624), .B(n11141), .Y(n2335) );
  NOR2X1TS U2717 ( .A(n10978), .B(n10276), .Y(n2917) );
  AOI211X1TS U2716 ( .A0(n9943), .A1(n11099), .B0(n2335), .C0(n2917), .Y(n3197) );
  OAI211X1TS U2715 ( .A0(n12474), .A1(n11901), .B0(n3196), .C0(n3197), .Y(
        n3195) );
  NOR2X1TS U2606 ( .A(n11632), .B(n10981), .Y(n2906) );
  OAI22X1TS U2604 ( .A0(n2895), .A1(n11625), .B0(n12174), .B1(n11484), .Y(
        n3151) );
  NOR2X1TS U2676 ( .A(n12146), .B(n11942), .Y(n1868) );
  OAI22X1TS U1959 ( .A0(n12482), .A1(n12477), .B0(n10978), .B1(n12353), .Y(
        n2680) );
  NOR2X1TS U2221 ( .A(n11899), .B(n2329), .Y(n2083) );
  NOR2X1TS U1729 ( .A(n11141), .B(n11905), .Y(n2088) );
  NOR2X1TS U1714 ( .A(n11582), .B(n9072), .Y(n2089) );
  NOR2X1TS U3126 ( .A(n10360), .B(n10363), .Y(n2668) );
  NOR2X1TS U3142 ( .A(n3306), .B(n2652), .Y(n2167) );
  NOR2X1TS U2343 ( .A(n10508), .B(n11526), .Y(n2639) );
  INVX2TS U3156 ( .A(n2765), .Y(n3316) );
  OAI22X1TS U1919 ( .A0(n11446), .A1(n12316), .B0(n10191), .B1(n11549), .Y(
        n2640) );
  AOI211X1TS U1918 ( .A0(n9956), .A1(n11816), .B0(n2639), .C0(n2640), .Y(n2632) );
  NOR2X1TS U3045 ( .A(n11561), .B(n10588), .Y(n2636) );
  NOR2X1TS U2385 ( .A(n11024), .B(n10949), .Y(n2637) );
  AOI21X1TS U1916 ( .A0(n11011), .A1(n11024), .B0(n2635), .Y(n2633) );
  INVX2TS U3084 ( .A(n9685), .Y(n2508) );
  NOR2X1TS U3078 ( .A(n11834), .B(n10596), .Y(n2160) );
  INVX2TS U3088 ( .A(n12339), .Y(n2510) );
  AOI22X1TS U3015 ( .A0(n1986), .A1(n11010), .B0(n11023), .B1(n9688), .Y(n3276) );
  NOR2X1TS U3023 ( .A(n11827), .B(n9956), .Y(n2776) );
  NOR2X1TS U3012 ( .A(n10619), .B(n12097), .Y(n3051) );
  AOI21X1TS U3011 ( .A0(n10630), .A1(n10510), .B0(n11063), .Y(n3280) );
  NOR2X1TS U3132 ( .A(n12623), .B(n11560), .Y(n2750) );
  OAI22X1TS U2037 ( .A0(n2750), .A1(n11835), .B0(n10187), .B1(n10624), .Y(
        n2047) );
  NOR2X1TS U3056 ( .A(n11062), .B(n10187), .Y(n3042) );
  NOR2X1TS U3052 ( .A(n1991), .B(n10191), .Y(n3027) );
  NOR2X1TS U2335 ( .A(n12341), .B(n10184), .Y(n2663) );
  NOR2X1TS U1939 ( .A(n11040), .B(n12288), .Y(n2059) );
  AOI22X1TS U1934 ( .A0(n11029), .A1(n12112), .B0(n10950), .B1(n10227), .Y(
        n2662) );
  OAI31X1TS U1933 ( .A0(n11526), .A1(n2660), .A2(n2661), .B0(n2662), .Y(n2659)
         );
  AOI211X1TS U1932 ( .A0(n12311), .A1(n12338), .B0(n2658), .C0(n2659), .Y(
        n2473) );
  NOR2X1TS U3139 ( .A(n11816), .B(n10223), .Y(n2777) );
  NOR2X1TS U2988 ( .A(n2777), .B(n10631), .Y(n2487) );
  INVX2TS U3044 ( .A(n2636), .Y(n2494) );
  AOI22X1TS U1810 ( .A0(n11561), .A1(n2491), .B0(n10224), .B1(n2159), .Y(n2490) );
  AOI211X1TS U1808 ( .A0(n11067), .A1(n2055), .B0(n2487), .C0(n2488), .Y(n2474) );
  NOR2X1TS U3027 ( .A(n10509), .B(n10191), .Y(n1980) );
  OAI22X1TS U3022 ( .A0(n2057), .A1(n11851), .B0(n2776), .B1(n11064), .Y(n3284) );
  AOI211X1TS U3021 ( .A0(n12615), .A1(n10516), .B0(n1980), .C0(n3284), .Y(
        n3281) );
  NOR2X1TS U3019 ( .A(n12112), .B(n10587), .Y(n2140) );
  OAI22X1TS U3018 ( .A0(n11834), .A1(n11016), .B0(n10962), .B1(n2140), .Y(
        n3283) );
  OAI211X1TS U3016 ( .A0(n11532), .A1(n11549), .B0(n3281), .C0(n3282), .Y(
        n2476) );
  INVX2TS U2471 ( .A(n9063), .Y(n2557) );
  NOR2X1TS U2530 ( .A(n2035), .B(n9844), .Y(n3001) );
  NOR2X1TS U2459 ( .A(n11005), .B(n12333), .Y(n1807) );
  NOR2X1TS U2576 ( .A(n2035), .B(n3139), .Y(n2194) );
  NOR2X1TS U2574 ( .A(n3002), .B(n12679), .Y(n2586) );
  OAI31X1TS U2456 ( .A0(n10584), .A1(n12092), .A2(n12323), .B0(n12188), .Y(
        n3114) );
  OAI31X1TS U2452 ( .A0(n10171), .A1(n11514), .A2(n10610), .B0(n12092), .Y(
        n3118) );
  AOI211X1TS U2450 ( .A0(n11057), .A1(n11424), .B0(n3116), .C0(n3117), .Y(
        n3115) );
  NOR2X1TS U2306 ( .A(n12323), .B(n11595), .Y(n2014) );
  OAI22X1TS U1573 ( .A0(n10606), .A1(n11589), .B0(n12565), .B1(n10685), .Y(
        n2024) );
  OAI22X1TS U1572 ( .A0(n2038), .A1(n12159), .B0(n11047), .B1(n9960), .Y(n2025) );
  AOI22X1TS U1571 ( .A0(n12360), .A1(n10679), .B0(n12333), .B1(n1806), .Y(
        n2037) );
  AOI22X1TS U1569 ( .A0(n12092), .A1(n11052), .B0(n10232), .B1(n11917), .Y(
        n2031) );
  NOR2X1TS U2447 ( .A(n10603), .B(n10011), .Y(n2974) );
  NOR2X1TS U2445 ( .A(n12332), .B(n11157), .Y(n2533) );
  AOI211X1TS U2440 ( .A0(n11512), .A1(n11955), .B0(n2974), .C0(n3109), .Y(
        n3108) );
  OAI211X1TS U2438 ( .A0(n10015), .A1(n10607), .B0(n3108), .C0(n2991), .Y(
        n2591) );
  NOR2X1TS U1905 ( .A(n12193), .B(n11911), .Y(n1804) );
  AOI211X1TS U1900 ( .A0(n10232), .A1(n11051), .B0(n2615), .C0(n2616), .Y(
        n2613) );
  OAI211X1TS U1899 ( .A0(n1804), .A1(n9968), .B0(n2613), .C0(n2614), .Y(n2592)
         );
  AOI22X1TS U1898 ( .A0(n2563), .A1(n12188), .B0(n11502), .B1(n11158), .Y(
        n2608) );
  NOR2X1TS U2248 ( .A(n10349), .B(n9055), .Y(n2612) );
  AOI22X1TS U1897 ( .A0(n2611), .A1(n2612), .B0(n10172), .B1(n9749), .Y(n2609)
         );
  INVX2TS U2245 ( .A(n9086), .Y(n2534) );
  NOR2X1TS U2308 ( .A(n11004), .B(n11519), .Y(n2607) );
  OAI22X1TS U1894 ( .A0(n2534), .A1(n12557), .B0(n2607), .B1(n11644), .Y(n2601) );
  OAI22X1TS U1892 ( .A0(n1824), .A1(n10291), .B0(n9995), .B1(n12159), .Y(n2603) );
  AOI22X1TS U1891 ( .A0(n12091), .A1(n10615), .B0(n12331), .B1(n11917), .Y(
        n2605) );
  OAI211X1TS U1890 ( .A0(n11590), .A1(n9959), .B0(n2605), .C0(n2606), .Y(n2604) );
  NOR2X1TS U2566 ( .A(n12565), .B(n11045), .Y(n2523) );
  NOR2X1TS U2546 ( .A(n11636), .B(n9928), .Y(n2995) );
  NOR2X1TS U2542 ( .A(n11948), .B(n10606), .Y(n3012) );
  AOI211X1TS U2541 ( .A0(n12093), .A1(n3000), .B0(n2995), .C0(n3012), .Y(n3141) );
  OAI211X1TS U2534 ( .A0(n10304), .A1(n11589), .B0(n3141), .C0(n3009), .Y(
        n3140) );
  AOI211X1TS U2533 ( .A0(n10611), .A1(n10180), .B0(n2523), .C0(n3140), .Y(
        n2595) );
  NOR2X1TS U2235 ( .A(n9996), .B(n10016), .Y(n2600) );
  NOR2X1TS U2416 ( .A(n12556), .B(n10694), .Y(n2994) );
  NOR2X1TS U2415 ( .A(n11636), .B(n9701), .Y(n2199) );
  AOI211X1TS U2414 ( .A0(n12333), .A1(n11506), .B0(n2994), .C0(n2199), .Y(
        n3091) );
  AOI211X1TS U2405 ( .A0(n12188), .A1(n12195), .B0(n3093), .C0(n3094), .Y(
        n3092) );
  NOR2X1TS U2386 ( .A(n10967), .B(n11042), .Y(n3035) );
  OAI22X1TS U2384 ( .A0(n2637), .A1(n10961), .B0(n9924), .B1(n11073), .Y(n3076) );
  AOI31X1TS U2381 ( .A0(sa03[6]), .A1(n10519), .A2(n9684), .B0(n3072), .Y(
        n3070) );
  OAI211X1TS U2380 ( .A0(n12118), .A1(n10620), .B0(n3070), .C0(n3071), .Y(
        n2751) );
  AOI22X1TS U2328 ( .A0(n11544), .A1(n11828), .B0(n12289), .B1(n11011), .Y(
        n3029) );
  OAI22X1TS U2059 ( .A0(n10960), .A1(n11017), .B0(n11080), .B1(n12118), .Y(
        n2772) );
  OAI22X1TS U2057 ( .A0(n11063), .A1(n11549), .B0(n11858), .B1(n12098), .Y(
        n2774) );
  OAI211X1TS U2053 ( .A0(n10961), .A1(n10598), .B0(n2770), .C0(n2771), .Y(
        n1953) );
  NOR2X1TS U2992 ( .A(n11458), .B(n12117), .Y(n2767) );
  NOR2X1TS U3003 ( .A(n12614), .B(n10224), .Y(n2769) );
  AOI211X1TS U2050 ( .A0(n10223), .A1(n12105), .B0(n2767), .C0(n2768), .Y(
        n2755) );
  AOI21X1TS U3114 ( .A0(n11081), .A1(n11550), .B0(n11524), .Y(n2759) );
  NOR2X1TS U3149 ( .A(n11009), .B(n10228), .Y(n2761) );
  NOR2X1TS U3001 ( .A(n12622), .B(n9955), .Y(n2153) );
  AOI211X1TS U2041 ( .A0(n9688), .A1(n2630), .B0(n2759), .C0(n2760), .Y(n2756)
         );
  OAI31X1TS U2040 ( .A0(n12111), .A1(n11562), .A2(n9094), .B0(n10228), .Y(
        n2757) );
  OAI22X1TS U1631 ( .A0(n11016), .A1(n11525), .B0(n11857), .B1(n12117), .Y(
        n2169) );
  AOI22X1TS U1629 ( .A0(n11041), .A1(n11030), .B0(n11023), .B1(n2058), .Y(
        n2165) );
  AOI211X1TS U1627 ( .A0(n11030), .A1(n2159), .B0(n2160), .C0(n2161), .Y(n2157) );
  OAI22X1TS U1625 ( .A0(n2140), .A1(n12318), .B0(n2153), .B1(n11036), .Y(n2152) );
  AOI211X1TS U1624 ( .A0(n11536), .A1(n2151), .B0(n1984), .C0(n2152), .Y(n2134) );
  AOI21X1TS U2356 ( .A0(n12309), .A1(n2628), .B0(n3051), .Y(n3049) );
  OAI211X1TS U2351 ( .A0(n10592), .A1(n11554), .B0(n2648), .C0(n3048), .Y(
        n3045) );
  OAI21X1TS U2349 ( .A0(n10966), .A1(n10183), .B0(n2061), .Y(n3047) );
  OAI211X1TS U2348 ( .A0(n12315), .A1(n11859), .B0(n2511), .C0(n3047), .Y(
        n3046) );
  NOR3X1TS U2347 ( .A(n3044), .B(n3045), .C(n3046), .Y(n2136) );
  AOI22X1TS U2394 ( .A0(n12340), .A1(n12614), .B0(n10520), .B1(n9094), .Y(
        n3077) );
  OAI31X1TS U2391 ( .A0(n10520), .A1(n12309), .A2(n11010), .B0(n10514), .Y(
        n3082) );
  NOR2X1TS U3006 ( .A(n12104), .B(n11561), .Y(n2149) );
  OAI22X1TS U1623 ( .A0(n2149), .A1(n10625), .B0(n2059), .B1(n12317), .Y(n2138) );
  NOR2X1TS U1912 ( .A(n10509), .B(n12116), .Y(n2146) );
  NOR4BX1TS U1619 ( .AN(n2136), .B(n2137), .C(n2138), .D(n2139), .Y(n2135) );
  INVX2TS U1555 ( .A(n1436), .Y(n1439) );
  NOR2X1TS U2071 ( .A(n10235), .B(n11524), .Y(n2782) );
  AOI31X1TS U2070 ( .A0(n11448), .A1(n10596), .A2(n11550), .B0(n2056), .Y(
        n2783) );
  OAI211X1TS U2068 ( .A0(n11079), .A1(n11852), .B0(n2791), .C0(n2512), .Y(
        n2784) );
  AOI22X1TS U2067 ( .A0(n12339), .A1(n11537), .B0(n12112), .B1(n2470), .Y(
        n2786) );
  OAI211X1TS U2064 ( .A0(n11460), .A1(n11530), .B0(n2786), .C0(n2787), .Y(
        n2785) );
  OAI22X1TS U1546 ( .A0(n11550), .A1(n12117), .B0(n1991), .B1(n11064), .Y(
        n1983) );
  OAI22X1TS U1545 ( .A0(n11555), .A1(n12098), .B0(n11851), .B1(n10619), .Y(
        n1985) );
  NOR3X1TS U1544 ( .A(n1983), .B(n1984), .C(n1985), .Y(n1977) );
  OAI32X1TS U1543 ( .A0(n1989), .A1(n1980), .A2(n12623), .B0(n11069), .B1(
        n1980), .Y(n1978) );
  OAI211X1TS U1542 ( .A0(n10236), .A1(n10626), .B0(n1977), .C0(n1978), .Y(
        n1954) );
  AOI21X1TS U1541 ( .A0(n10631), .A1(n11857), .B0(n11075), .Y(n1962) );
  NOR2X1TS U2379 ( .A(n11441), .B(n11537), .Y(n1964) );
  AOI22X1TS U3106 ( .A0(n10515), .A1(n9689), .B0(n9955), .B1(n10228), .Y(n1967) );
  AOI22X1TS U2376 ( .A0(n11029), .A1(n11827), .B0(n12615), .B1(n10183), .Y(
        n3067) );
  OAI211X1TS U2375 ( .A0(n1964), .A1(n11016), .B0(n3066), .C0(n3067), .Y(n3052) );
  OAI211X1TS U2373 ( .A0(n12317), .A1(n9924), .B0(n3065), .C0(n2634), .Y(n3059) );
  AOI211X1TS U2367 ( .A0(n12622), .A1(n10223), .B0(n3059), .C0(n3060), .Y(
        n2742) );
  AOI211X1TS U2361 ( .A0(n9956), .A1(n2491), .B0(n2487), .C0(n3057), .Y(n3056)
         );
  NOR4BX1TS U1536 ( .AN(n1952), .B(n1953), .C(n1954), .D(n1955), .Y(n1312) );
  AOI31X1TS U1535 ( .A0(n12166), .A1(n10662), .A2(n2293), .B0(n11572), .Y(
        n1889) );
  NOR2X1TS U2793 ( .A(n10247), .B(n1939), .Y(n1951) );
  OAI22X1TS U1534 ( .A0(n9108), .A1(n11865), .B0(n1951), .B1(n12458), .Y(n1890) );
  AOI22X1TS U1532 ( .A0(n10239), .A1(n11085), .B0(n9975), .B1(n1927), .Y(n1940) );
  OAI21X1TS U1531 ( .A0(n12126), .A1(n10637), .B0(n11871), .Y(n1941) );
  OAI211X1TS U1530 ( .A0(n1757), .A1(n10244), .B0(n1940), .C0(n1941), .Y(n1891) );
  NOR2X1TS U2839 ( .A(n12346), .B(n11612), .Y(n2827) );
  NOR2X1TS U2022 ( .A(n11601), .B(n11428), .Y(n2294) );
  OAI22X1TS U1698 ( .A0(n11608), .A1(n12086), .B0(n11881), .B1(n1925), .Y(
        n2295) );
  AOI211X1TS U1697 ( .A0(n10578), .A1(n10561), .B0(n2294), .C0(n2295), .Y(
        n2283) );
  OAI21X1TS U1696 ( .A0(n10575), .A1(n12085), .B0(n2292), .Y(n2290) );
  AOI211X1TS U1695 ( .A0(n10260), .A1(n11116), .B0(n2289), .C0(n2290), .Y(
        n2284) );
  OAI21X1TS U1693 ( .A0(n11881), .A1(n12167), .B0(n2288), .Y(n2287) );
  AOI211X1TS U1692 ( .A0(n11931), .A1(n1740), .B0(n2114), .C0(n2287), .Y(n2285) );
  AOI22X1TS U1528 ( .A0(n11089), .A1(n1937), .B0(n1908), .B1(n1762), .Y(n1913)
         );
  AOI22X1TS U1527 ( .A0(n12133), .A1(n1933), .B0(n11095), .B1(n1935), .Y(n1914) );
  AOI211X1TS U1525 ( .A0(n9741), .A1(n1927), .B0(n1929), .C0(n1930), .Y(n1915)
         );
  NOR2X1TS U2840 ( .A(n12468), .B(n11865), .Y(n1918) );
  NOR2X1TS U2808 ( .A(n12123), .B(n12301), .Y(n2805) );
  AOI211X1TS U2079 ( .A0(n9724), .A1(n10564), .B0(n2730), .C0(n2804), .Y(n2802) );
  AOI22X1TS U1523 ( .A0(n12605), .A1(n11567), .B0(n10247), .B1(n1927), .Y(
        n1924) );
  NOR3X1TS U1519 ( .A(n1910), .B(n1911), .C(n1912), .Y(n1732) );
  AOI21X1TS U2902 ( .A0(n11120), .A1(n10252), .B0(n10641), .Y(n2860) );
  OAI211X1TS U2141 ( .A0(n12466), .A1(n10641), .B0(n2862), .C0(n2863), .Y(
        n2861) );
  AOI211X1TS U2140 ( .A0(n12302), .A1(n1937), .B0(n2860), .C0(n2861), .Y(n2859) );
  OAI211X1TS U2139 ( .A0(n10654), .A1(n11429), .B0(n2858), .C0(n2859), .Y(
        n2857) );
  AOI211X1TS U2138 ( .A0(n10988), .A1(n9976), .B0(n2109), .C0(n2857), .Y(n1893) );
  AOI22X1TS U1687 ( .A0(n9740), .A1(n10987), .B0(n10247), .B1(n10295), .Y(
        n2276) );
  AOI211X1TS U1680 ( .A0(n12124), .A1(n9947), .B0(n2264), .C0(n2265), .Y(n1894) );
  NOR2X1TS U2023 ( .A(n11863), .B(n10252), .Y(n1897) );
  OAI211X1TS U2095 ( .A0(n11120), .A1(n10658), .B0(n2816), .C0(n2817), .Y(
        n1898) );
  NOR4BX1TS U1515 ( .AN(n1896), .B(n1897), .C(n1898), .D(n1899), .Y(n1895) );
  AOI31X1TS U1511 ( .A0(n12173), .A1(n10675), .A2(n11149), .B0(n11583), .Y(
        n1826) );
  NOR2X1TS U2596 ( .A(n10271), .B(n12296), .Y(n1888) );
  OAI22X1TS U1510 ( .A0(n9112), .A1(n11888), .B0(n1888), .B1(n12475), .Y(n1827) );
  AOI22X1TS U1508 ( .A0(n10263), .A1(n11099), .B0(n9987), .B1(n1864), .Y(n1877) );
  OAI21X1TS U1507 ( .A0(n12140), .A1(n10645), .B0(n11894), .Y(n1878) );
  OAI211X1TS U1506 ( .A0(n1719), .A1(n10268), .B0(n1877), .C0(n1878), .Y(n1828) );
  AOI22X1TS U2181 ( .A0(n9631), .A1(n11152), .B0(n11847), .B1(n2686), .Y(n2900) );
  NOR2X1TS U2642 ( .A(n12353), .B(n11631), .Y(n2903) );
  AOI211X1TS U2179 ( .A0(n10528), .A1(n12372), .B0(n2903), .C0(n2904), .Y(
        n2901) );
  NOR2X1TS U1980 ( .A(n11619), .B(n11434), .Y(n2361) );
  OAI22X1TS U1733 ( .A0(n11626), .A1(n12079), .B0(n11906), .B1(n1862), .Y(
        n2362) );
  AOI211X1TS U1732 ( .A0(n10552), .A1(n10534), .B0(n2361), .C0(n2362), .Y(
        n2350) );
  OAI21X1TS U1731 ( .A0(n10548), .A1(n12078), .B0(n2359), .Y(n2357) );
  AOI211X1TS U1730 ( .A0(n10283), .A1(n11137), .B0(n2356), .C0(n2357), .Y(
        n2351) );
  OAI21X1TS U1728 ( .A0(n11907), .A1(n12173), .B0(n2355), .Y(n2354) );
  AOI211X1TS U1727 ( .A0(n11943), .A1(n10539), .B0(n2088), .C0(n2354), .Y(
        n2352) );
  AOI22X1TS U1504 ( .A0(n11105), .A1(n1874), .B0(n11110), .B1(n1724), .Y(n1850) );
  AOI22X1TS U1503 ( .A0(n12144), .A1(n1870), .B0(n11111), .B1(n1872), .Y(n1851) );
  AOI211X1TS U1501 ( .A0(n9745), .A1(n1864), .B0(n1866), .C0(n1867), .Y(n1852)
         );
  NOR2X1TS U2643 ( .A(n12484), .B(n11889), .Y(n1855) );
  NOR2X1TS U2611 ( .A(n12137), .B(n12295), .Y(n2881) );
  AOI211X1TS U2154 ( .A0(n9728), .A1(n10538), .B0(n2697), .C0(n2880), .Y(n2878) );
  NOR3X1TS U1495 ( .A(n1847), .B(n1848), .C(n1849), .Y(n1694) );
  AOI21X1TS U2705 ( .A0(n11143), .A1(n10276), .B0(n10650), .Y(n2936) );
  OAI21X1TS U2217 ( .A0(n10534), .A1(n12295), .B0(n11895), .Y(n2938) );
  OAI211X1TS U2216 ( .A0(n12482), .A1(n10650), .B0(n2938), .C0(n2939), .Y(
        n2937) );
  AOI211X1TS U2215 ( .A0(n1876), .A1(n1874), .B0(n2936), .C0(n2937), .Y(n2935)
         );
  OAI211X1TS U2214 ( .A0(n10666), .A1(n11435), .B0(n2934), .C0(n2935), .Y(
        n2933) );
  AOI211X1TS U2213 ( .A0(n10972), .A1(n9988), .B0(n2083), .C0(n2933), .Y(n1830) );
  AOI211X1TS U1715 ( .A0(n12140), .A1(n9943), .B0(n2331), .C0(n2332), .Y(n1831) );
  NOR2X1TS U1981 ( .A(n11889), .B(n10275), .Y(n1834) );
  OAI211X1TS U2170 ( .A0(n11142), .A1(n10671), .B0(n2892), .C0(n2893), .Y(
        n1835) );
  NOR4BX1TS U1491 ( .AN(n1833), .B(n1834), .C(n1835), .D(n1836), .Y(n1832) );
  NOR4X1TS U1489 ( .A(n1826), .B(n1827), .C(n1828), .D(n1829), .Y(n1417) );
  NOR2X1TS U2277 ( .A(n11047), .B(n9959), .Y(n2979) );
  AOI22X1TS U2271 ( .A0(n11821), .A1(n10168), .B0(n12358), .B1(n2984), .Y(
        n2983) );
  OAI22X1TS U1834 ( .A0(n2533), .A1(n11643), .B0(n2534), .B1(n2540), .Y(n2524)
         );
  NOR2X1TS U2527 ( .A(n11423), .B(n11594), .Y(n2531) );
  AOI22X1TS U1832 ( .A0(n12360), .A1(n12153), .B0(n12331), .B1(n10611), .Y(
        n2527) );
  NOR2X1TS U2500 ( .A(n10693), .B(n10175), .Y(n2529) );
  NOR2X1TS U1875 ( .A(n10176), .B(n10303), .Y(n2530) );
  AOI211X1TS U1831 ( .A0(n11003), .A1(n11500), .B0(n2529), .C0(n2530), .Y(
        n2528) );
  OAI211X1TS U1830 ( .A0(n11636), .A1(n9963), .B0(n2527), .C0(n2528), .Y(n2526) );
  AOI22X1TS U2301 ( .A0(n1693), .A1(n12091), .B0(n12152), .B1(n11954), .Y(
        n3003) );
  AOI22X1TS U2300 ( .A0(n12154), .A1(n12332), .B0(n12194), .B1(n10611), .Y(
        n3004) );
  OAI22X1TS U1881 ( .A0(n2038), .A1(n11047), .B0(n10007), .B1(n10685), .Y(
        n1795) );
  NOR2X1TS U2504 ( .A(n10007), .B(n10602), .Y(n2992) );
  AOI21X1TS U2278 ( .A0(n10615), .A1(n2185), .B0(n2987), .Y(n2203) );
  AOI21X1TS U1856 ( .A0(n11947), .A1(n11644), .B0(n9996), .Y(n2550) );
  OAI211X1TS U1851 ( .A0(n2552), .A1(n11948), .B0(n2553), .C0(n2554), .Y(n2551) );
  AOI211X1TS U1850 ( .A0(n1803), .A1(n1802), .B0(n2550), .C0(n2551), .Y(n2204)
         );
  NOR2X1TS U2464 ( .A(n2587), .B(n9700), .Y(n2214) );
  AOI21X1TS U1846 ( .A0(n9051), .A1(n10088), .B0(n11919), .Y(n2216) );
  AOI211X1TS U1653 ( .A0(n12187), .A1(n2213), .B0(n2214), .C0(n2215), .Y(n2205) );
  OAI211X1TS U2302 ( .A0(n10694), .A1(n11638), .B0(n3010), .C0(n3011), .Y(
        n2207) );
  INVX2TS U1477 ( .A(n9254), .Y(n1338) );
  INVX2TS U3328 ( .A(n3396), .Y(n3395) );
  AOI22X1TS U5677 ( .A0(n9954), .A1(n10146), .B0(n11207), .B1(n10497), .Y(
        n6164) );
  NOR2X1TS U5676 ( .A(n5298), .B(n11674), .Y(n5410) );
  NOR2X1TS U5672 ( .A(n9287), .B(n6040), .Y(n5780) );
  AOI211X1TS U5670 ( .A0(n10555), .A1(n6187), .B0(n5780), .C0(n6188), .Y(n6184) );
  AOI211X1TS U5658 ( .A0(n11685), .A1(n11335), .B0(n6175), .C0(n6176), .Y(
        n6172) );
  NOR2X1TS U5568 ( .A(n9954), .B(n9998), .Y(n5416) );
  NOR2X1TS U5558 ( .A(n6039), .B(n10185), .Y(n5611) );
  OAI22X1TS U5406 ( .A0(n5746), .A1(n12019), .B0(n5769), .B1(n10974), .Y(n5768) );
  NOR4BX1TS U5405 ( .AN(n5765), .B(n5766), .C(n5767), .D(n5768), .Y(n5734) );
  AOI22X1TS U5830 ( .A0(n11718), .A1(n10249), .B0(n10968), .B1(n10478), .Y(
        n6354) );
  NOR2X1TS U5829 ( .A(n11347), .B(n10182), .Y(n5668) );
  OAI31X1TS U5810 ( .A0(n9407), .A1(n11999), .A2(n11742), .B0(n10941), .Y(
        n6356) );
  NOR2X1TS U5782 ( .A(n10969), .B(n10576), .Y(n5676) );
  OAI22X1TS U5404 ( .A0(n5763), .A1(n5994), .B0(n5676), .B1(n5657), .Y(n5738)
         );
  AOI22X1TS U5395 ( .A0(n11353), .A1(n12536), .B0(n11329), .B1(n10479), .Y(
        n5741) );
  AOI22X1TS U5394 ( .A0(n10969), .A1(n9977), .B0(n5760), .B1(n11741), .Y(n5742) );
  OAI211X1TS U5391 ( .A0(n5660), .A1(n9723), .B0(n5734), .C0(n5735), .Y(n1776)
         );
  AOI22X1TS U5171 ( .A0(n5203), .A1(n9259), .B0(n12673), .B1(n5206), .Y(n5250)
         );
  OAI21X1TS U5432 ( .A0(n12210), .A1(n10522), .B0(n5822), .Y(n5771) );
  OAI32X1TS U5431 ( .A0(n10043), .A1(n10154), .A2(n9985), .B0(n10824), .B1(
        n10190), .Y(n5816) );
  OAI22X1TS U5560 ( .A0(n10417), .A1(n5309), .B0(n12441), .B1(n5630), .Y(n6031) );
  AOI22X1TS U5430 ( .A0(n11685), .A1(n10146), .B0(n11228), .B1(n11979), .Y(
        n5818) );
  OAI211X1TS U5426 ( .A0(n5809), .A1(n12497), .B0(n5810), .C0(n5811), .Y(n5773) );
  OAI211X1TS U5563 ( .A0(n6043), .A1(n10990), .B0(n6044), .C0(n6045), .Y(n6042) );
  AOI211X1TS U5562 ( .A0(n10562), .A1(n10246), .B0(n6041), .C0(n6042), .Y(
        n6038) );
  OAI211X1TS U5561 ( .A0(n5416), .A1(n6040), .B0(n6037), .C0(n6038), .Y(n5788)
         );
  AOI211X1TS U5423 ( .A0(n10491), .A1(n5803), .B0(n5804), .C0(n5805), .Y(n5801) );
  AOI211X1TS U5411 ( .A0(n11378), .A1(n5779), .B0(n5780), .C0(n5781), .Y(n5777) );
  AOI22X1TS U5879 ( .A0(n10582), .A1(n5692), .B0(n11688), .B1(n6426), .Y(n6396) );
  OAI22X1TS U5875 ( .A0(n6388), .A1(n11251), .B0(n9715), .B1(n12417), .Y(n6072) );
  OAI211X1TS U5853 ( .A0(n5494), .A1(n9360), .B0(n6402), .C0(n6403), .Y(n6401)
         );
  NOR4BX1TS U5852 ( .AN(n6399), .B(n5467), .C(n6400), .D(n6401), .Y(n6398) );
  OAI22X1TS U5460 ( .A0(n5864), .A1(n10210), .B0(n5865), .B1(n10214), .Y(n5846) );
  NOR2X1TS U5713 ( .A(n10909), .B(n11270), .Y(n5696) );
  AOI22X1TS U5450 ( .A0(n10864), .A1(n11270), .B0(n10994), .B1(n11002), .Y(
        n5850) );
  OAI211X1TS U5437 ( .A0(n9715), .A1(n12025), .B0(n5826), .C0(n5827), .Y(n1621) );
  INVX2TS U5436 ( .A(n1621), .Y(n1619) );
  AOI21X1TS U5725 ( .A0(n9384), .A1(n9533), .B0(n11222), .Y(n6134) );
  AOI211X1TS U5624 ( .A0(n11698), .A1(n12589), .B0(n5509), .C0(n6137), .Y(
        n6136) );
  NOR2X1TS U5749 ( .A(n10937), .B(n11318), .Y(n5721) );
  OAI22X1TS U5747 ( .A0(n5721), .A1(n12424), .B0(n5387), .B1(n10511), .Y(n6258) );
  AOI22X1TS U5745 ( .A0(n12248), .A1(n11971), .B0(n11325), .B1(n11014), .Y(
        n6266) );
  AOI22X1TS U5743 ( .A0(n12519), .A1(n9961), .B0(n11013), .B1(n9734), .Y(n6263) );
  OAI211X1TS U5742 ( .A0(n6262), .A1(n11366), .B0(n6263), .C0(n6264), .Y(n6261) );
  AOI22X1TS U5621 ( .A0(n12048), .A1(n9308), .B0(n9961), .B1(n9372), .Y(n6127)
         );
  NOR2X1TS U5620 ( .A(n12589), .B(n11971), .Y(n5723) );
  AOI211X1TS U5617 ( .A0(n9633), .A1(n9734), .B0(n6129), .C0(n6130), .Y(n6128)
         );
  NOR4BX1TS U5615 ( .AN(n6121), .B(n6122), .C(n6123), .D(n6124), .Y(n5709) );
  OAI211X1TS U5613 ( .A0(n11390), .A1(n10470), .B0(n6120), .C0(n5898), .Y(
        n6095) );
  OAI22X1TS U5950 ( .A0(n6460), .A1(n11299), .B0(n9719), .B1(n12425), .Y(n6116) );
  OAI22X1TS U5734 ( .A0(n11215), .A1(n12402), .B0(n9707), .B1(n11390), .Y(
        n6243) );
  OAI21X1TS U5732 ( .A0(n12250), .A1(n11006), .B0(n11012), .Y(n6248) );
  OAI211X1TS U5730 ( .A0(n12400), .A1(n10920), .B0(n6248), .C0(n5519), .Y(
        n6245) );
  NOR4BX1TS U5600 ( .AN(n5709), .B(n6095), .C(n6096), .D(n6097), .Y(n1574) );
  OAI22X1TS U5164 ( .A0(n5248), .A1(n12748), .B0(n12685), .B1(n5249), .Y(N180)
         );
  AOI22X1TS U5653 ( .A0(n10145), .A1(n6162), .B0(n11981), .B1(n5783), .Y(n6145) );
  OAI22X1TS U5640 ( .A0(n5632), .A1(n5616), .B0(n10149), .B1(n10959), .Y(n5406) );
  NOR3X1TS U5634 ( .A(n6142), .B(n5605), .C(n6143), .Y(n1531) );
  AOI211X1TS U5797 ( .A0(n10250), .A1(n5995), .B0(n5563), .C0(n6336), .Y(n6328) );
  AOI22X1TS U5796 ( .A0(n12061), .A1(n6335), .B0(n5573), .B1(n12544), .Y(n5664) );
  OAI22X1TS U5794 ( .A0(n12020), .A1(n9388), .B0(n12013), .B1(n12007), .Y(
        n6332) );
  NOR3X1TS U5790 ( .A(n6326), .B(n5737), .C(n6327), .Y(n1648) );
  INVX2TS U5631 ( .A(n5226), .Y(n5225) );
  AOI22X1TS U5196 ( .A0(n5225), .A1(n9260), .B0(n12673), .B1(n5226), .Y(n5266)
         );
  AOI22X1TS U5842 ( .A0(n12583), .A1(n10886), .B0(n11275), .B1(n9297), .Y(
        n5695) );
  NOR4BX1TS U5838 ( .AN(n5695), .B(n6385), .C(n6386), .D(n6387), .Y(n6380) );
  NOR4BX1TS U5833 ( .AN(n5430), .B(n5468), .C(n5845), .D(n6379), .Y(n1612) );
  INVX2TS U5832 ( .A(n1612), .Y(n1614) );
  OAI22X1TS U5189 ( .A0(n5264), .A1(n12746), .B0(n12685), .B1(n5265), .Y(N177)
         );
  AOI22X1TS U3948 ( .A0(n12566), .A1(n10460), .B0(n10875), .B1(n10134), .Y(
        n4549) );
  AOI211X1TS U3942 ( .A0(n10802), .A1(n9691), .B0(n4576), .C0(n4577), .Y(n4574) );
  OAI31X1TS U3928 ( .A0(n11701), .A1(n10806), .A2(n4536), .B0(n9687), .Y(n4551) );
  AOI211X1TS U3915 ( .A0(n11702), .A1(n4532), .B0(n4533), .C0(n4534), .Y(n4527) );
  OAI22X1TS U3914 ( .A0(n3953), .A1(n10770), .B0(n10783), .B1(n10144), .Y(
        n3906) );
  NOR3X1TS U3908 ( .A(n4524), .B(n3938), .C(n4525), .Y(n1781) );
  INVX2TS U3748 ( .A(n3429), .Y(n3428) );
  AOI22X1TS U3316 ( .A0(n3428), .A1(n9074), .B0(n12674), .B1(n3429), .Y(n3468)
         );
  OAI22X1TS U3308 ( .A0(n3466), .A1(n12751), .B0(n12688), .B1(n3467), .Y(N241)
         );
  AOI22X1TS U3290 ( .A0(n3406), .A1(n9073), .B0(n12674), .B1(n3409), .Y(n3452)
         );
  AOI211X1TS U3547 ( .A0(n10433), .A1(n4017), .B0(n4018), .C0(n4019), .Y(n4015) );
  OAI21X1TS U3539 ( .A0(n9929), .A1(n10787), .B0(n4002), .Y(n3994) );
  OAI211X1TS U3536 ( .A0(n12276), .A1(n3821), .B0(n3997), .C0(n3998), .Y(n3995) );
  AOI211X1TS U3535 ( .A0(n11799), .A1(n10156), .B0(n3994), .C0(n3995), .Y(
        n3971) );
  OAI211X1TS U3530 ( .A0(n3985), .A1(n11709), .B0(n3987), .C0(n3988), .Y(n3975) );
  INVX2TS U3524 ( .A(n9191), .Y(n3365) );
  AOI22X1TS U3288 ( .A0(n3365), .A1(n9316), .B0(n9314), .B1(n9191), .Y(n3454)
         );
  OAI22X1TS U3577 ( .A0(n4064), .A1(n10106), .B0(n4065), .B1(n10110), .Y(n4046) );
  AOI22X1TS U3567 ( .A0(n10906), .A1(n11333), .B0(n10760), .B1(n10768), .Y(
        n4050) );
  OAI211X1TS U3554 ( .A0(n9659), .A1(n12008), .B0(n4026), .C0(n4027), .Y(n1635) );
  INVX2TS U3553 ( .A(n1635), .Y(n1633) );
  AOI22X1TS U3673 ( .A0(n11987), .A1(n9115), .B0(n9910), .B1(n9165), .Y(n4217)
         );
  NOR2X1TS U3672 ( .A(n12580), .B(n12053), .Y(n3893) );
  NOR4BX1TS U3667 ( .AN(n4211), .B(n4212), .C(n4213), .D(n4214), .Y(n3879) );
  OAI211X1TS U3665 ( .A0(n11237), .A1(n10438), .B0(n4210), .C0(n4098), .Y(
        n4185) );
  NOR4BX1TS U3652 ( .AN(n3879), .B(n4185), .C(n4186), .D(n4187), .Y(n1588) );
  OAI22X1TS U3283 ( .A0(n3450), .A1(n12751), .B0(n12688), .B1(n3451), .Y(N244)
         );
  OAI22X1TS U3743 ( .A0(n9678), .A1(n12022), .B0(n9640), .B1(n3665), .Y(n4329)
         );
  AOI22X1TS U3736 ( .A0(n11703), .A1(n4324), .B0(n3672), .B1(n3911), .Y(n4323)
         );
  AOI211X1TS U3727 ( .A0(n10460), .A1(n4300), .B0(n4301), .C0(n4302), .Y(n4299) );
  OAI211X1TS U3726 ( .A0(n4297), .A1(n12208), .B0(n4298), .C0(n4299), .Y(n4288) );
  NOR4BX1TS U3720 ( .AN(n4286), .B(n4287), .C(n4288), .D(n4289), .Y(n3904) );
  INVX2TS U3718 ( .A(n1787), .Y(n1785) );
  AOI22X1TS U3300 ( .A0(n9073), .A1(n3415), .B0(n3416), .B1(n12674), .Y(n3458)
         );
  AOI211X1TS U3648 ( .A0(n11749), .A1(n12585), .B0(n3688), .C0(n4183), .Y(
        n4182) );
  AOI22X1TS U3645 ( .A0(n12001), .A1(n9107), .B0(n9905), .B1(n9158), .Y(n4173)
         );
  NOR2X1TS U3644 ( .A(n9636), .B(n12057), .Y(n3868) );
  AOI211X1TS U3641 ( .A0(n9636), .A1(n9646), .B0(n4175), .C0(n4176), .Y(n4174)
         );
  NOR4BX1TS U3639 ( .AN(n4167), .B(n4168), .C(n4169), .D(n4170), .Y(n3854) );
  OAI211X1TS U3637 ( .A0(n11243), .A1(n10447), .B0(n4166), .C0(n4042), .Y(
        n4141) );
  NOR4BX1TS U3624 ( .AN(n3854), .B(n4141), .C(n4142), .D(n4143), .Y(n1630) );
  OAI22X1TS U3292 ( .A0(n3456), .A1(n12751), .B0(n12688), .B1(n3457), .Y(N243)
         );
  AOI21X1TS U5769 ( .A0(n10722), .A1(n9392), .B0(n10946), .Y(n5991) );
  AOI22X1TS U5531 ( .A0(n10550), .A1(n5995), .B0(n10940), .B1(n9352), .Y(n5992) );
  OAI211X1TS U5529 ( .A0(n5991), .A1(n11372), .B0(n5992), .C0(n5993), .Y(n5990) );
  AOI211X1TS U5528 ( .A0(n11997), .A1(n5988), .B0(n5989), .C0(n5990), .Y(n5975) );
  OAI211X1TS U5777 ( .A0(n6311), .A1(n10233), .B0(n6312), .C0(n6313), .Y(n6310) );
  OAI211X1TS U5775 ( .A0(n5676), .A1(n5578), .B0(n6307), .C0(n6308), .Y(n5979)
         );
  AOI22X1TS U5527 ( .A0(n12544), .A1(n10178), .B0(n10238), .B1(n12535), .Y(
        n5986) );
  AOI22X1TS U5525 ( .A0(n10545), .A1(n10193), .B0(n12434), .B1(n10479), .Y(
        n5982) );
  AOI32X1TS U5524 ( .A0(n5982), .A1(n10234), .A2(n9727), .B0(n12006), .B1(
        n5982), .Y(n5981) );
  OAI211X1TS U5518 ( .A0(n11989), .A1(n9727), .B0(n5969), .C0(n5970), .Y(n5968) );
  OAI21X1TS U5768 ( .A0(n11753), .A1(n11747), .B0(n6301), .Y(n6300) );
  AOI211X1TS U5767 ( .A0(n10545), .A1(n11717), .B0(n6299), .C0(n6300), .Y(
        n5946) );
  AOI211X1TS U5511 ( .A0(n10940), .A1(n5955), .B0(n5956), .C0(n5957), .Y(n5947) );
  AOI22X1TS U5774 ( .A0(n12054), .A1(n11998), .B0(n11354), .B1(n10478), .Y(
        n6303) );
  OAI211X1TS U5770 ( .A0(n5668), .A1(n5984), .B0(n6303), .C0(n6304), .Y(n5951)
         );
  AOI22X1TS U5181 ( .A0(n9259), .A1(n5212), .B0(n5213), .B1(n12673), .Y(n5256)
         );
  OAI22X1TS U5553 ( .A0(n12442), .A1(n10500), .B0(n12212), .B1(n10957), .Y(
        n6017) );
  AOI22X1TS U5550 ( .A0(n10558), .A1(n9994), .B0(n11378), .B1(n10242), .Y(
        n6022) );
  OAI22X1TS U5547 ( .A0(n6014), .A1(n10825), .B0(n9312), .B1(n11402), .Y(n6001) );
  AOI211X1TS U5539 ( .A0(n11342), .A1(n9284), .B0(n6001), .C0(n6002), .Y(n5999) );
  NOR3X1TS U5536 ( .A(n5788), .B(n5997), .C(n5998), .Y(n5166) );
  OAI22X1TS U5740 ( .A0(n10571), .A1(n9707), .B0(n10470), .B1(n11313), .Y(
        n6250) );
  OAI22X1TS U5739 ( .A0(n5543), .A1(n10541), .B0(n11289), .B1(n12399), .Y(
        n6251) );
  AOI211X1TS U5737 ( .A0(n10439), .A1(n11319), .B0(n6255), .C0(n6256), .Y(
        n6254) );
  OAI211X1TS U5736 ( .A0(n10166), .A1(n10218), .B0(n6253), .C0(n6254), .Y(
        n6252) );
  AOI31X1TS U5726 ( .A0(n9303), .A1(n11215), .A2(n10873), .B0(n5514), .Y(n6231) );
  OAI22X1TS U5724 ( .A0(n9302), .A1(n9775), .B0(n6134), .B1(n11301), .Y(n6233)
         );
  AOI22X1TS U5723 ( .A0(n12243), .A1(n10912), .B0(n11293), .B1(n9371), .Y(
        n6236) );
  OAI211X1TS U5717 ( .A0(n6235), .A1(n5557), .B0(n6236), .C0(n6237), .Y(n6234)
         );
  AOI21X1TS U5689 ( .A0(n9380), .A1(n9326), .B0(n11211), .Y(n6090) );
  AOI211X1TS U5596 ( .A0(n11680), .A1(n12581), .B0(n5443), .C0(n6093), .Y(
        n6092) );
  OAI22X1TS U5711 ( .A0(n5696), .A1(n12416), .B0(n5348), .B1(n10505), .Y(n6218) );
  AOI22X1TS U5709 ( .A0(n12225), .A1(n11974), .B0(n11277), .B1(n11002), .Y(
        n6226) );
  AOI22X1TS U5707 ( .A0(n12503), .A1(n9957), .B0(n11001), .B1(n9730), .Y(n6223) );
  OAI211X1TS U5706 ( .A0(n6222), .A1(n11360), .B0(n6223), .C0(n6224), .Y(n6221) );
  AOI22X1TS U5593 ( .A0(n12035), .A1(n9298), .B0(n9957), .B1(n9363), .Y(n6083)
         );
  NOR2X1TS U5592 ( .A(n12582), .B(n11974), .Y(n5698) );
  AOI211X1TS U5589 ( .A0(n9635), .A1(n9731), .B0(n6085), .C0(n6086), .Y(n6084)
         );
  NOR4BX1TS U5587 ( .AN(n6077), .B(n6078), .C(n6079), .D(n6080), .Y(n5684) );
  OAI211X1TS U5585 ( .A0(n11384), .A1(n6384), .B0(n6076), .C0(n5842), .Y(n6051) );
  OAI22X1TS U5698 ( .A0(n11203), .A1(n12386), .B0(n9703), .B1(n11384), .Y(
        n6203) );
  OAI22X1TS U5697 ( .A0(n11360), .A1(n10858), .B0(n10568), .B1(n10507), .Y(
        n6204) );
  OAI21X1TS U5696 ( .A0(n12227), .A1(n10994), .B0(n11000), .Y(n6208) );
  NOR4BX1TS U5572 ( .AN(n5684), .B(n6051), .C(n6052), .D(n6053), .Y(n1616) );
  OAI22X1TS U5173 ( .A0(n5254), .A1(n12747), .B0(n12685), .B1(n5255), .Y(N179)
         );
  INVX2TS U4186 ( .A(n9126), .Y(n4023) );
  AOI22X1TS U3680 ( .A0(n4023), .A1(n3421), .B0(n3422), .B1(n9125), .Y(n4229)
         );
  OAI22X1TS U3619 ( .A0(n4137), .A1(n12750), .B0(n12687), .B1(n4138), .Y(N227)
         );
  OAI22X1TS U3499 ( .A0(n9921), .A1(n12573), .B0(n9639), .B1(n12381), .Y(n3899) );
  OAI211X1TS U3496 ( .A0(n3919), .A1(n9650), .B0(n3921), .C0(n3922), .Y(n3900)
         );
  AOI31X1TS U3489 ( .A0(n9654), .A1(n3896), .A2(n10420), .B0(n10815), .Y(n3873) );
  OAI22X1TS U3487 ( .A0(n3892), .A1(n10809), .B0(n3893), .B1(n11255), .Y(n3874) );
  AOI32X1TS U3486 ( .A0(n3889), .A1(n3890), .A2(n3891), .B0(n11297), .B1(n3890), .Y(n3875) );
  AOI22X1TS U3483 ( .A0(n10901), .A1(n3887), .B0(n10804), .B1(n12237), .Y(
        n3885) );
  AOI211X1TS U3481 ( .A0(n11285), .A1(n10889), .B0(n3881), .C0(n3882), .Y(
        n3880) );
  AOI31X1TS U7174 ( .A0(n9491), .A1(n11522), .A2(n11528), .B0(n11868), .Y(
        n7302) );
  OAI22X1TS U7173 ( .A0(n7333), .A1(n10661), .B0(n9492), .B1(n11109), .Y(n7323) );
  AOI22X1TS U7172 ( .A0(n11517), .A1(n7330), .B0(n11861), .B1(n7332), .Y(n7327) );
  OAI211X1TS U7171 ( .A0(n10030), .A1(n11103), .B0(n7327), .C0(n7328), .Y(
        n7324) );
  OAI211X1TS U7169 ( .A0(n7317), .A1(n11510), .B0(n7319), .C0(n7320), .Y(n7303) );
  OAI22X1TS U7168 ( .A0(n10286), .A1(n10647), .B0(n10652), .B1(n10657), .Y(
        n7312) );
  AOI211X1TS U7167 ( .A0(n10281), .A1(n11096), .B0(n7311), .C0(n7312), .Y(
        n7308) );
  NOR4BX1TS U7165 ( .AN(n7301), .B(n7302), .C(n7303), .D(n7304), .Y(n6965) );
  OAI22X1TS U3211 ( .A0(n3373), .A1(n12752), .B0(n12689), .B1(n3374), .Y(N273)
         );
  AOI22X1TS U3203 ( .A0(n3365), .A1(n9338), .B0(n9336), .B1(n9192), .Y(n3361)
         );
  OAI22X1TS U3198 ( .A0(n3357), .A1(n12752), .B0(n12690), .B1(n3358), .Y(N275)
         );
  AOI31X1TS U5383 ( .A0(n9718), .A1(n5726), .A2(n10513), .B0(n10923), .Y(n5703) );
  OAI22X1TS U5381 ( .A0(n5722), .A1(n10930), .B0(n5723), .B1(n11367), .Y(n5704) );
  AOI22X1TS U5917 ( .A0(n12589), .A1(n10914), .B0(n11323), .B1(n9307), .Y(
        n5720) );
  AOI32X1TS U5380 ( .A0(n5719), .A1(n5720), .A2(n5721), .B0(n11307), .B1(n5720), .Y(n5705) );
  AOI211X1TS U5375 ( .A0(n11317), .A1(n10879), .B0(n5711), .C0(n5712), .Y(
        n5710) );
  AOI31X1TS U5371 ( .A0(n9714), .A1(n5701), .A2(n10507), .B0(n10896), .Y(n5678) );
  OAI22X1TS U5369 ( .A0(n5697), .A1(n10904), .B0(n5698), .B1(n11359), .Y(n5679) );
  AOI32X1TS U5368 ( .A0(n5694), .A1(n5695), .A2(n5696), .B0(n11257), .B1(n5695), .Y(n5680) );
  OAI22X1TS U5704 ( .A0(n10566), .A1(n9703), .B0(n10462), .B1(n11265), .Y(
        n6210) );
  OAI22X1TS U5703 ( .A0(n5477), .A1(n10530), .B0(n11241), .B1(n12383), .Y(
        n6211) );
  AOI211X1TS U5701 ( .A0(n10421), .A1(n11271), .B0(n6215), .C0(n6216), .Y(
        n6214) );
  OAI211X1TS U5700 ( .A0(n10158), .A1(n10210), .B0(n6213), .C0(n6214), .Y(
        n6212) );
  AOI211X1TS U5363 ( .A0(n11269), .A1(n10864), .B0(n5686), .C0(n5687), .Y(
        n5685) );
  OAI22X1TS U5761 ( .A0(n10483), .A1(n10198), .B0(n11018), .B1(n10230), .Y(
        n6280) );
  AOI22X1TS U5760 ( .A0(n10970), .A1(n9973), .B0(n10549), .B1(n10201), .Y(
        n6282) );
  AOI22X1TS U5758 ( .A0(n11724), .A1(n6286), .B0(n5574), .B1(n10250), .Y(n6284) );
  NOR4BX1TS U5756 ( .AN(n6278), .B(n6279), .C(n6280), .D(n6281), .Y(n5650) );
  AOI22X1TS U1146 ( .A0(n1305), .A1(n1303), .B0(n1304), .B1(n9779), .Y(n1301)
         );
  NOR2X1TS U2612 ( .A(n10553), .B(n11488), .Y(n2920) );
  AOI211X1TS U2195 ( .A0(n12138), .A1(n10300), .B0(n2917), .C0(n2918), .Y(
        n2883) );
  AOI21X1TS U2700 ( .A0(n10276), .A1(n12352), .B0(n11434), .Y(n2915) );
  NOR2X1TS U2609 ( .A(n10283), .B(n10203), .Y(n2313) );
  AOI211X1TS U2193 ( .A0(n11941), .A1(n9745), .B0(n2915), .C0(n2916), .Y(n2884) );
  AOI22X1TS U2168 ( .A0(n10973), .A1(n2100), .B0(n11936), .B1(n2890), .Y(n2396) );
  OAI31X1TS U2165 ( .A0(n1702), .A1(n12296), .A2(n9761), .B0(n1845), .Y(n2889)
         );
  NOR4BX1TS U2163 ( .AN(n1695), .B(n1847), .C(n1835), .D(n2886), .Y(n2885) );
  OAI22X1TS U1725 ( .A0(n12484), .A1(n10671), .B0(n12173), .B1(n10212), .Y(
        n2348) );
  AOI21X1TS U1724 ( .A0(n11895), .A1(n2100), .B0(n2348), .Y(n2347) );
  OAI31X1TS U1723 ( .A0(n9713), .A1(n2346), .A2(n2087), .B0(n2347), .Y(n2299)
         );
  NOR2X1TS U1750 ( .A(n11477), .B(n10982), .Y(n2315) );
  OAI22X1TS U1713 ( .A0(n12175), .A1(n12476), .B0(n12352), .B1(n10544), .Y(
        n2316) );
  NOR2X1TS U2674 ( .A(n9631), .B(n9943), .Y(n2327) );
  NOR2X1TS U1964 ( .A(n10676), .B(n10671), .Y(n2322) );
  OAI32X1TS U1709 ( .A0(n11936), .A1(n2322), .A2(n11153), .B0(n9943), .B1(
        n2322), .Y(n2321) );
  OAI211X1TS U1708 ( .A0(n10208), .A1(n9072), .B0(n2320), .C0(n2321), .Y(n2317) );
  NOR2X1TS U1952 ( .A(n11887), .B(n10268), .Y(n2309) );
  OAI22X1TS U1706 ( .A0(n2311), .A1(n1882), .B0(n2313), .B1(n10212), .Y(n2310)
         );
  AOI211X1TS U1705 ( .A0(n11894), .A1(n11106), .B0(n2309), .C0(n2310), .Y(
        n2301) );
  NOR2X1TS U2622 ( .A(n11583), .B(n12353), .Y(n2304) );
  AOI211X1TS U1703 ( .A0(n10553), .A1(n1720), .B0(n2304), .C0(n2305), .Y(n2302) );
  OAI22X1TS U3610 ( .A0(n4120), .A1(n10114), .B0(n4121), .B1(n10118), .Y(n4102) );
  AOI22X1TS U3600 ( .A0(n10887), .A1(n11284), .B0(n10772), .B1(n10778), .Y(
        n4106) );
  OAI211X1TS U3587 ( .A0(n9655), .A1(n11993), .B0(n4082), .C0(n4083), .Y(n1593) );
  INVX2TS U3586 ( .A(n1593), .Y(n1591) );
  INVX2TS U3551 ( .A(n3355), .Y(n3354) );
  AOI211X1TS U3372 ( .A0(n10932), .A1(n3601), .B0(n3602), .C0(n3603), .Y(n3346) );
  OAI22X1TS U3254 ( .A0(n3423), .A1(n12751), .B0(n12689), .B1(n3424), .Y(N257)
         );
  AOI22X1TS U5123 ( .A0(n5203), .A1(n12664), .B0(n5205), .B1(n5206), .Y(n5200)
         );
  AOI22X1TS U5954 ( .A0(n5511), .A1(n5717), .B0(n11706), .B1(n6498), .Y(n6468)
         );
  OAI211X1TS U5928 ( .A0(n5560), .A1(n9368), .B0(n6474), .C0(n6475), .Y(n6473)
         );
  NOR4BX1TS U5927 ( .AN(n6471), .B(n5533), .C(n6472), .D(n6473), .Y(n6470) );
  OAI22X1TS U5493 ( .A0(n5920), .A1(n10218), .B0(n5921), .B1(n10222), .Y(n5902) );
  OAI211X1TS U5470 ( .A0(n9719), .A1(n12040), .B0(n5882), .C0(n5883), .Y(n1579) );
  INVX2TS U5469 ( .A(n1579), .Y(n1577) );
  OAI22X1TS U5117 ( .A0(n5198), .A1(n12758), .B0(n12686), .B1(n5199), .Y(N196)
         );
  NOR4BX1TS U5913 ( .AN(n5720), .B(n6457), .C(n6458), .D(n6459), .Y(n6452) );
  NOR4BX1TS U5908 ( .AN(n5496), .B(n5534), .C(n5901), .D(n6451), .Y(n1570) );
  OAI22X1TS U5136 ( .A0(n5220), .A1(n12749), .B0(n12686), .B1(n5221), .Y(N193)
         );
  OAI22X1TS U3236 ( .A0(n3401), .A1(n12752), .B0(n12689), .B1(n3402), .Y(N260)
         );
  INVX2TS U5135 ( .A(n5177), .Y(n5176) );
  AOI22X1TS U5099 ( .A0(n9267), .A1(n5176), .B0(n5177), .B1(n12675), .Y(n5170)
         );
  OAI22X1TS U5091 ( .A0(n5168), .A1(n12758), .B0(n12686), .B1(n5169), .Y(N209)
         );
  INVX2TS U5434 ( .A(n5149), .Y(n5148) );
  AOI22X1TS U5075 ( .A0(n9268), .A1(n5148), .B0(n5149), .B1(n12675), .Y(n5143)
         );
  OAI22X1TS U5068 ( .A0(n5141), .A1(n12750), .B0(n12687), .B1(n5142), .Y(N212)
         );
  AOI22X1TS U1877 ( .A0(n11823), .A1(n12181), .B0(n12326), .B1(n2228), .Y(
        n2580) );
  NOR2X1TS U1876 ( .A(n10693), .B(n11642), .Y(n2195) );
  AOI211X1TS U1874 ( .A0(n10680), .A1(n12331), .B0(n2195), .C0(n2530), .Y(
        n2581) );
  AOI211X1TS U1871 ( .A0(n11507), .A1(n11003), .B0(n2578), .C0(n2579), .Y(
        n1655) );
  AOI22X1TS U2478 ( .A0(n11501), .A1(n12093), .B0(n12151), .B1(n10583), .Y(
        n3124) );
  AOI21X1TS U2475 ( .A0(n11508), .A1(n11422), .B0(n3121), .Y(n2568) );
  NOR2X1TS U2508 ( .A(n2611), .B(n12180), .Y(n1670) );
  AOI211X1TS U2460 ( .A0(n11004), .A1(n2221), .B0(n2214), .C0(n3119), .Y(n3102) );
  NOR2X1TS U2426 ( .A(n12152), .B(n11500), .Y(n1672) );
  INVX2TS U1425 ( .A(n9261), .Y(n1325) );
  INVX2TS U1423 ( .A(n1418), .Y(n1419) );
  AOI22X1TS U1203 ( .A0(n1417), .A1(n1418), .B0(n1419), .B1(n1420), .Y(n1416)
         );
  OAI22X1TS U3243 ( .A0(n3410), .A1(n12752), .B0(n12689), .B1(n3411), .Y(N259)
         );
  AOI31X1TS U5690 ( .A0(n9293), .A1(n11203), .A2(n10857), .B0(n12028), .Y(
        n6191) );
  OAI22X1TS U5688 ( .A0(n9292), .A1(n9771), .B0(n6090), .B1(n11253), .Y(n6193)
         );
  AOI22X1TS U5687 ( .A0(n12220), .A1(n10884), .B0(n11245), .B1(n9363), .Y(
        n6196) );
  OAI211X1TS U5681 ( .A0(n6195), .A1(n5491), .B0(n6196), .C0(n6197), .Y(n6194)
         );
  AOI22X1TS U6987 ( .A0(n9456), .A1(n1297), .B0(n1298), .B1(n12678), .Y(n6968)
         );
  OAI22X1TS U6979 ( .A0(n6966), .A1(n12740), .B0(n12683), .B1(n6967), .Y(N145)
         );
  AOI22X1TS U6972 ( .A0(n9455), .A1(n1277), .B0(n1278), .B1(n12678), .Y(n6956)
         );
  OAI22X1TS U6964 ( .A0(n6954), .A1(n12741), .B0(n12684), .B1(n6955), .Y(N147)
         );
  AOI22X1TS U6963 ( .A0(n9455), .A1(n6951), .B0(n6952), .B1(n12678), .Y(n6946)
         );
  OAI22X1TS U6956 ( .A0(n6944), .A1(n12742), .B0(n12684), .B1(n6945), .Y(N148)
         );
  NOR2X1TS U3007 ( .A(n10948), .B(n10184), .Y(n3043) );
  AOI21X1TS U2344 ( .A0(n11555), .A1(n11447), .B0(n11035), .Y(n3038) );
  OAI211X1TS U2340 ( .A0(n11853), .A1(n11017), .B0(n3040), .C0(n3041), .Y(
        n3039) );
  AOI31X1TS U2336 ( .A0(n11852), .A1(n11064), .A2(n2781), .B0(n11556), .Y(
        n3020) );
  OAI211X1TS U2331 ( .A0(n2663), .A1(n11525), .B0(n3033), .C0(n3034), .Y(n3021) );
  OAI211X1TS U2320 ( .A0(n11524), .A1(n11081), .B0(n2509), .C0(n3023), .Y(
        n3022) );
  INVX2TS U2317 ( .A(n1413), .Y(n1412) );
  NOR2X1TS U2812 ( .A(n11132), .B(n10637), .Y(n2856) );
  AOI22X1TS U2134 ( .A0(n1939), .A1(n10296), .B0(n11869), .B1(n2252), .Y(n2852) );
  OAI22X1TS U2133 ( .A0(n10993), .A1(n10998), .B0(n12087), .B1(n11882), .Y(
        n2855) );
  AOI211X1TS U2132 ( .A0(n9740), .A1(n12602), .B0(n2854), .C0(n2855), .Y(n2853) );
  AOI22X1TS U1460 ( .A0(n11117), .A1(n9757), .B0(n11925), .B1(n1768), .Y(n1759) );
  OAI211X1TS U1458 ( .A0(n1757), .A1(n10653), .B0(n1759), .C0(n1760), .Y(n1736) );
  OAI22X1TS U1457 ( .A0(n12166), .A1(n1754), .B0(n2293), .B1(n10658), .Y(n1737) );
  OAI22X1TS U1456 ( .A0(n12468), .A1(n11606), .B0(n11600), .B1(n12460), .Y(
        n1738) );
  NOR2X1TS U2874 ( .A(n10663), .B(n11464), .Y(n1748) );
  NOR2X1TS U1777 ( .A(n11465), .B(n10999), .Y(n2248) );
  OAI22X1TS U1678 ( .A0(n12168), .A1(n12459), .B0(n12348), .B1(n10570), .Y(
        n2249) );
  NOR2X1TS U2871 ( .A(n9627), .B(n9947), .Y(n2260) );
  NOR2X1TS U2006 ( .A(n10662), .B(n10658), .Y(n2255) );
  OAI32X1TS U1674 ( .A0(n11925), .A1(n2255), .A2(n11131), .B0(n9948), .B1(
        n2255), .Y(n2254) );
  OAI211X1TS U1673 ( .A0(n10215), .A1(n9079), .B0(n2253), .C0(n2254), .Y(n2250) );
  INVX2TS U1451 ( .A(n9265), .Y(n1315) );
  INVX2TS U1449 ( .A(n9776), .Y(n1358) );
  AOI22X1TS U1240 ( .A0(n1358), .A1(n1325), .B0(n9262), .B1(n9776), .Y(n1478)
         );
  NOR2X1TS U2525 ( .A(n11912), .B(n11157), .Y(n2961) );
  OAI22X1TS U2524 ( .A0(n2531), .A1(n11590), .B0(n2961), .B1(n11948), .Y(n3131) );
  AOI21X1TS U2515 ( .A0(n9932), .A1(n10288), .B0(n12556), .Y(n3133) );
  AOI211X1TS U2499 ( .A0(n12181), .A1(n10179), .B0(n2992), .C0(n2529), .Y(
        n3136) );
  OAI211X1TS U2498 ( .A0(n9721), .A1(n12161), .B0(n3135), .C0(n3136), .Y(n3134) );
  NOR2X1TS U2493 ( .A(n11637), .B(n2220), .Y(n2975) );
  OAI22X1TS U2491 ( .A0(n12557), .A1(n1669), .B0(n10176), .B1(n10011), .Y(
        n3129) );
  AOI211X1TS U2490 ( .A0(n11913), .A1(n10003), .B0(n2975), .C0(n3129), .Y(
        n3083) );
  AOI211X1TS U2422 ( .A0(n11057), .A1(n2577), .B0(n3098), .C0(n2615), .Y(n3096) );
  OAI211X1TS U2398 ( .A0(n1809), .A1(n9967), .B0(n3087), .C0(n3088), .Y(n3086)
         );
  INVX2TS U2395 ( .A(n9227), .Y(n1480) );
  AOI22X1TS U3197 ( .A0(n12676), .A1(n3354), .B0(n3355), .B1(n9080), .Y(n3349)
         );
  OAI22X1TS U3190 ( .A0(n3347), .A1(n12753), .B0(n12690), .B1(n3348), .Y(N276)
         );
  AOI22X1TS U2905 ( .A0(n10635), .A1(n2453), .B0(n10987), .B1(n1933), .Y(n3226) );
  AOI21X1TS U2897 ( .A0(n10252), .A1(n12348), .B0(n11428), .Y(n2839) );
  OAI22X1TS U2870 ( .A0(n1931), .A1(n10654), .B0(n2260), .B1(n12346), .Y(n3243) );
  OAI211X1TS U2867 ( .A0(n10220), .A1(n12085), .B0(n3242), .C0(n2867), .Y(
        n2414) );
  AOI22X1TS U2863 ( .A0(n12605), .A1(n10636), .B0(n12133), .B1(n12303), .Y(
        n3240) );
  NOR2X1TS U2819 ( .A(n11572), .B(n1947), .Y(n2237) );
  AOI211X1TS U2816 ( .A0(n12131), .A1(n10260), .B0(n2237), .C0(n3219), .Y(
        n3218) );
  AOI32X1TS U2815 ( .A0(n12168), .A1(n3218), .A2(n12466), .B0(n10641), .B1(
        n3218), .Y(n3202) );
  NOR2X1TS U2811 ( .A(n11090), .B(n2252), .Y(n2436) );
  OAI22X1TS U2810 ( .A0(n2856), .A1(n10574), .B0(n2436), .B1(n10219), .Y(n3215) );
  NOR2X1TS U2809 ( .A(n10580), .B(n11496), .Y(n2844) );
  NOR2X1TS U2806 ( .A(n10259), .B(n10200), .Y(n2246) );
  OAI22X1TS U2794 ( .A0(n11571), .A1(n12087), .B0(n11122), .B1(n11471), .Y(
        n3208) );
  AOI211X1TS U2791 ( .A0(n9971), .A1(n2734), .B0(n3208), .C0(n3209), .Y(n2437)
         );
  AOI22X1TS U2789 ( .A0(n12604), .A1(n11130), .B0(n11871), .B1(n11925), .Y(
        n3207) );
  OAI211X1TS U2787 ( .A0(n10640), .A1(n11602), .B0(n3207), .C0(n2288), .Y(
        n2434) );
  AOI211X1TS U2786 ( .A0(n12123), .A1(n11116), .B0(n3206), .C0(n2434), .Y(
        n3205) );
  NOR2X1TS U2615 ( .A(n11154), .B(n10645), .Y(n2932) );
  AOI22X1TS U2209 ( .A0(n12295), .A1(n10299), .B0(n11893), .B1(n11578), .Y(
        n2928) );
  OAI22X1TS U2208 ( .A0(n10977), .A1(n1880), .B0(n12078), .B1(n11906), .Y(
        n2931) );
  AOI211X1TS U2207 ( .A0(n9744), .A1(n12599), .B0(n2930), .C0(n2931), .Y(n2929) );
  AOI22X1TS U1447 ( .A0(n11137), .A1(n9760), .B0(n11935), .B1(n1730), .Y(n1721) );
  OAI211X1TS U1445 ( .A0(n1719), .A1(n10667), .B0(n1721), .C0(n1722), .Y(n1698) );
  OAI22X1TS U1444 ( .A0(n12175), .A1(n1716), .B0(n11148), .B1(n10671), .Y(
        n1699) );
  OAI22X1TS U1443 ( .A0(n12485), .A1(n11624), .B0(n11618), .B1(n12474), .Y(
        n1700) );
  NOR2X1TS U2677 ( .A(n10675), .B(n11476), .Y(n1710) );
  INVX2TS U1438 ( .A(n9230), .Y(n1475) );
  OAI22X1TS U1311 ( .A0(n9228), .A1(n9231), .B0(n1475), .B1(n1480), .Y(n1317)
         );
  AOI22X1TS U3130 ( .A0(n10967), .A1(n2514), .B0(n11069), .B1(n2159), .Y(n3286) );
  AOI211X1TS U3104 ( .A0(n10949), .A1(n3031), .B0(n2759), .C0(n3320), .Y(n3287) );
  AOI22X1TS U3100 ( .A0(n11817), .A1(n12111), .B0(n10950), .B1(n12308), .Y(
        n3317) );
  AOI22X1TS U3094 ( .A0(n11829), .A1(n10224), .B0(n12105), .B1(n11536), .Y(
        n3318) );
  OAI22X1TS U3080 ( .A0(n2499), .A1(n12316), .B0(n9105), .B1(n10523), .Y(n3290) );
  AOI211X1TS U3033 ( .A0(n10520), .A1(n2494), .B0(n3293), .C0(n2503), .Y(n3292) );
  NOR2X1TS U3004 ( .A(n12290), .B(n10588), .Y(n2465) );
  NOR2X1TS U2997 ( .A(n10596), .B(n11074), .Y(n2779) );
  AOI32X1TS U2994 ( .A0(n9692), .A1(n3271), .A2(n12099), .B0(n11017), .B1(
        n3271), .Y(n3270) );
  AOI211X1TS U2993 ( .A0(n10227), .A1(n12110), .B0(n2779), .C0(n3270), .Y(
        n2501) );
  AOI211X1TS U2989 ( .A0(n12622), .A1(n11815), .B0(n2767), .C0(n3269), .Y(
        n3264) );
  OAI211X1TS U2984 ( .A0(n12097), .A1(n10188), .B0(n3268), .C0(n3074), .Y(
        n2462) );
  OAI22X1TS U2983 ( .A0(n9104), .A1(n11525), .B0(n9692), .B1(n11857), .Y(n3267) );
  OAI22X1TS U2287 ( .A0(n2531), .A1(n12161), .B0(n2617), .B1(n9960), .Y(n2970)
         );
  AOI22X1TS U2265 ( .A0(n10172), .A1(n12093), .B0(n11454), .B1(n11954), .Y(
        n2976) );
  AOI22X1TS U2264 ( .A0(n12333), .A1(n2549), .B0(n11518), .B1(n2978), .Y(n2977) );
  NOR4BX1TS U2258 ( .AN(n2968), .B(n2969), .C(n2970), .D(n2971), .Y(n2963) );
  AOI22X1TS U2257 ( .A0(n10171), .A1(n11157), .B0(n11500), .B1(n12323), .Y(
        n2966) );
  OAI22X1TS U2254 ( .A0(n10000), .A1(n9963), .B0(n11643), .B1(n10303), .Y(
        n2965) );
  OAI211X1TS U2252 ( .A0(n1662), .A1(n10956), .B0(n2963), .C0(n2964), .Y(n2519) );
  NOR4BX1TS U2241 ( .AN(n2957), .B(n2958), .C(n2959), .D(n2960), .Y(n2945) );
  AOI22X1TS U2238 ( .A0(n10168), .A1(n2561), .B0(n10231), .B1(n2619), .Y(n2956) );
  AOI211X1TS U2233 ( .A0(n11502), .A1(n11423), .B0(n2600), .C0(n2953), .Y(
        n2946) );
  OAI211X1TS U2231 ( .A0(n10693), .A1(n10004), .B0(n2950), .C0(n2951), .Y(
        n2226) );
  INVX2TS U2223 ( .A(n1472), .Y(n1471) );
  AOI22X1TS U5261 ( .A0(n9953), .A1(n11670), .B0(n11227), .B1(n11675), .Y(
        n5421) );
  AOI211X1TS U5254 ( .A0(n10834), .A1(n5399), .B0(n5400), .C0(n5401), .Y(n5140) );
  AOI22X1TS U4099 ( .A0(n4023), .A1(n3434), .B0(n3435), .B1(n9125), .Y(n4521)
         );
  OAI22X1TS U3901 ( .A0(n4519), .A1(n12750), .B0(n12687), .B1(n4520), .Y(N225)
         );
  OAI22X1TS U5766 ( .A0(n6297), .A1(n10226), .B0(n6298), .B1(n9981), .Y(n6291)
         );
  AOI22X1TS U5765 ( .A0(n12432), .A1(n6295), .B0(n12300), .B1(n9352), .Y(n6293) );
  OAI211X1TS U5764 ( .A0(n11982), .A1(n11989), .B0(n6293), .C0(n6294), .Y(
        n6292) );
  OAI211X1TS U5762 ( .A0(n5991), .A1(n12007), .B0(n5946), .C0(n6290), .Y(n6270) );
  AOI211X1TS U5753 ( .A0(n12542), .A1(n12055), .B0(n5569), .C0(n6275), .Y(
        n6273) );
  OAI31X1TS U5752 ( .A0(n10970), .A1(n11997), .A2(n5586), .B0(n12534), .Y(
        n6274) );
  AOI22X1TS U5134 ( .A0(n5217), .A1(n5218), .B0(n5219), .B1(n12658), .Y(n5216)
         );
  AOI22X1TS U2708 ( .A0(n2308), .A1(n2409), .B0(n10973), .B1(n1870), .Y(n3166)
         );
  OAI22X1TS U2673 ( .A0(n1868), .A1(n10667), .B0(n2327), .B1(n12352), .Y(n3183) );
  OAI211X1TS U2670 ( .A0(n10212), .A1(n12080), .B0(n3182), .C0(n2943), .Y(
        n2370) );
  AOI22X1TS U2666 ( .A0(n9632), .A1(n10645), .B0(n12144), .B1(n12297), .Y(
        n3180) );
  AOI211X1TS U2641 ( .A0(n1712), .A1(n9064), .B0(n1855), .C0(n2903), .Y(n3172)
         );
  OAI22X1TS U2597 ( .A0(n11582), .A1(n12080), .B0(n11142), .B1(n11483), .Y(
        n3148) );
  AOI211X1TS U2594 ( .A0(n9983), .A1(n2701), .B0(n3148), .C0(n3149), .Y(n2393)
         );
  AOI22X1TS U2592 ( .A0(n12601), .A1(n11153), .B0(n11895), .B1(n11936), .Y(
        n3147) );
  OAI211X1TS U2590 ( .A0(n10649), .A1(n11620), .B0(n3147), .C0(n2355), .Y(
        n2390) );
  OAI22X1TS U1235 ( .A0(n9230), .A1(n9266), .B0(n1315), .B1(n1475), .Y(n1437)
         );
  INVX2TS U1234 ( .A(n1437), .Y(n1438) );
  AOI22X1TS U1233 ( .A0(n1470), .A1(n1471), .B0(n1472), .B1(n1473), .Y(n1469)
         );
  AOI22X1TS U5066 ( .A0(n9263), .A1(n1774), .B0(n1776), .B1(n5139), .Y(n5137)
         );
  AOI22X1TS U1132 ( .A0(n12661), .A1(n1277), .B0(n1278), .B1(n1279), .Y(n1269)
         );
  OAI22X1TS U1127 ( .A0(n1266), .A1(n12757), .B0(n12682), .B1(n1268), .Y(N99)
         );
  AOI22X1TS U1258 ( .A0(n1436), .A1(n9269), .B0(n12672), .B1(n1439), .Y(n1493)
         );
  AOI211X1TS U2120 ( .A0(n12123), .A1(n10295), .B0(n2841), .C0(n2842), .Y(
        n2807) );
  AOI211X1TS U2118 ( .A0(n11930), .A1(n9741), .B0(n2839), .C0(n2840), .Y(n2808) );
  AOI22X1TS U2093 ( .A0(n10986), .A1(n2126), .B0(n11923), .B1(n2814), .Y(n2440) );
  OAI31X1TS U2090 ( .A0(n10565), .A1(n12301), .A2(n9756), .B0(n1908), .Y(n2813) );
  NOR4BX1TS U2088 ( .AN(n1733), .B(n1910), .C(n1898), .D(n2810), .Y(n2809) );
  OAI22X1TS U1690 ( .A0(n12467), .A1(n10659), .B0(n12169), .B1(n10220), .Y(
        n2281) );
  AOI21X1TS U1689 ( .A0(n11871), .A1(n2126), .B0(n2281), .Y(n2280) );
  OAI31X1TS U1688 ( .A0(n9717), .A1(n2279), .A2(n2113), .B0(n2280), .Y(n2232)
         );
  NOR2X1TS U1994 ( .A(n11865), .B(n10244), .Y(n2242) );
  OAI22X1TS U1671 ( .A0(n2244), .A1(n1945), .B0(n2246), .B1(n10220), .Y(n2243)
         );
  AOI211X1TS U1670 ( .A0(n11869), .A1(n11088), .B0(n2242), .C0(n2243), .Y(
        n2234) );
  AOI211X1TS U1668 ( .A0(n10580), .A1(n11084), .B0(n2237), .C0(n2238), .Y(
        n2235) );
  NOR4X1TS U1666 ( .A(n1911), .B(n2231), .C(n2232), .D(n2233), .Y(n1342) );
  INVX2TS U1665 ( .A(n1342), .Y(n1343) );
  OAI22X1TS U1963 ( .A0(n12174), .A1(n11477), .B0(n12483), .B1(n11436), .Y(
        n2689) );
  AOI211X1TS U1962 ( .A0(n1876), .A1(n11135), .B0(n2322), .C0(n2689), .Y(n2394) );
  AOI22X1TS U1754 ( .A0(n10538), .A1(n1874), .B0(n10300), .B1(n2096), .Y(n2373) );
  NOR3X1TS U1752 ( .A(n2389), .B(n2390), .C(n2391), .Y(n2374) );
  AOI211X1TS U1744 ( .A0(n10527), .A1(n9988), .B0(n2377), .C0(n2378), .Y(n2376) );
  NOR4X1TS U1742 ( .A(n2370), .B(n2075), .C(n2371), .D(n2372), .Y(n1445) );
  OAI21X1TS U1845 ( .A0(n12562), .A1(n11636), .B0(n2545), .Y(n2544) );
  AOI221X1TS U1844 ( .A0(n2563), .A1(n2559), .B0(n11058), .B1(n12323), .C0(
        n2544), .Y(n2182) );
  AOI21X1TS U1837 ( .A0(n12325), .A1(n11918), .B0(n2537), .Y(n2536) );
  INVX2TS U1635 ( .A(n9246), .Y(n1372) );
  INVX2TS U1741 ( .A(n1445), .Y(n1447) );
  OAI22X1TS U1252 ( .A0(n1491), .A1(n12754), .B0(n12691), .B1(n1492), .Y(N52)
         );
  OAI22X1TS U2005 ( .A0(n12167), .A1(n11464), .B0(n12469), .B1(n11430), .Y(
        n2722) );
  AOI211X1TS U2004 ( .A0(n12302), .A1(n11115), .B0(n2255), .C0(n2722), .Y(
        n2438) );
  AOI22X1TS U1781 ( .A0(n10564), .A1(n1937), .B0(n10296), .B1(n2122), .Y(n2417) );
  OAI22X1TS U1780 ( .A0(n2436), .A1(n10216), .B0(n10654), .B1(n12459), .Y(
        n2435) );
  NOR3X1TS U1779 ( .A(n2433), .B(n2434), .C(n2435), .Y(n2418) );
  AOI211X1TS U1771 ( .A0(n1750), .A1(n9975), .B0(n2421), .C0(n2422), .Y(n2420)
         );
  NOR4X1TS U1769 ( .A(n2414), .B(n2101), .C(n2415), .D(n2416), .Y(n1351) );
  INVX2TS U1768 ( .A(n1351), .Y(n1354) );
  OAI22X1TS U1208 ( .A0(n1428), .A1(n12760), .B0(n12694), .B1(n1429), .Y(N68)
         );
  OAI22X1TS U5076 ( .A0(n5151), .A1(n12758), .B0(n12687), .B1(n5152), .Y(N211)
         );
  AOI22X1TS U1157 ( .A0(n1325), .A1(n9616), .B0(n9614), .B1(n9261), .Y(n1324)
         );
  OAI22X1TS U1153 ( .A0(n1319), .A1(n12755), .B0(n12694), .B1(n1320), .Y(N86)
         );
  AOI22X1TS U5112 ( .A0(n5190), .A1(n5191), .B0(n5192), .B1(n9170), .Y(n5189)
         );
  AOI22X1TS U1245 ( .A0(n1338), .A1(n1418), .B0(n1419), .B1(n9255), .Y(n1484)
         );
  INVX2TS U6069 ( .A(n9318), .Y(n5823) );
  AOI22X1TS U5532 ( .A0(n5823), .A1(n5218), .B0(n5219), .B1(n9317), .Y(n5941)
         );
  OAI22X1TS U5502 ( .A0(n5937), .A1(n12744), .B0(n12684), .B1(n5938), .Y(N163)
         );
  AOI22X1TS U7100 ( .A0(n6927), .A1(n7008), .B0(n7007), .B1(n9794), .Y(n7096)
         );
  OAI22X1TS U7082 ( .A0(n7092), .A1(n12735), .B0(n12682), .B1(n7093), .Y(N115)
         );
  AOI22X1TS U3231 ( .A0(n3394), .A1(n3395), .B0(n3396), .B1(n9163), .Y(n3393)
         );
  AOI22X1TS U3277 ( .A0(n3346), .A1(n3395), .B0(n3396), .B1(n9187), .Y(n3444)
         );
  OAI22X1TS U2010 ( .A0(n2260), .A1(n9979), .B0(n2725), .B1(n11612), .Y(n2724)
         );
  AOI31X1TS U2008 ( .A0(n9109), .A1(n2286), .A2(n12468), .B0(n11471), .Y(n2704) );
  OAI211X1TS U2002 ( .A0(n2449), .A1(n10255), .B0(n2438), .C0(n2721), .Y(n2706) );
  AOI22X1TS U1986 ( .A0(n12604), .A1(n10260), .B0(n11929), .B1(n9976), .Y(
        n2709) );
  INVX2TS U1982 ( .A(n9251), .Y(n1369) );
  OAI22X1TS U1968 ( .A0(n2327), .A1(n9991), .B0(n2692), .B1(n11630), .Y(n2691)
         );
  AOI31X1TS U1966 ( .A0(n9113), .A1(n2353), .A2(n12484), .B0(n11483), .Y(n2671) );
  OAI211X1TS U1960 ( .A0(n2405), .A1(n10279), .B0(n2394), .C0(n2688), .Y(n2673) );
  AOI22X1TS U1944 ( .A0(n9631), .A1(n10284), .B0(n11942), .B1(n9987), .Y(n2676) );
  OAI22X1TS U1931 ( .A0(n2499), .A1(n11062), .B0(n9104), .B1(n11530), .Y(n2653) );
  AOI22X1TS U1930 ( .A0(n11817), .A1(n2494), .B0(n12104), .B1(n2657), .Y(n2656) );
  OAI211X1TS U1929 ( .A0(n9090), .A1(n11549), .B0(n2655), .C0(n2656), .Y(n2654) );
  AOI211X1TS U1928 ( .A0(n12339), .A1(n11009), .B0(n2653), .C0(n2654), .Y(
        n2620) );
  AOI31X1TS U1926 ( .A0(n11447), .A1(n9923), .A2(n9105), .B0(n11073), .Y(n2645) );
  OAI211X1TS U1924 ( .A0(n9693), .A1(n10510), .B0(n2647), .C0(n2648), .Y(n2496) );
  AOI211X1TS U1923 ( .A0(n10966), .A1(n2493), .B0(n2645), .C0(n2496), .Y(n2621) );
  OAI22X1TS U1922 ( .A0(n11034), .A1(n10188), .B0(n10621), .B1(n11532), .Y(
        n2644) );
  AOI221X1TS U1921 ( .A0(n11544), .A1(n10948), .B0(n11022), .B1(n11067), .C0(
        n2644), .Y(n2623) );
  OAI22X1TS U1911 ( .A0(n11015), .A1(n11531), .B0(n10620), .B1(n11526), .Y(
        n2627) );
  OAI211X1TS U1909 ( .A0(n2060), .A1(n10192), .B0(n2625), .C0(n2626), .Y(n2495) );
  NOR4BX1TS U1908 ( .AN(n2623), .B(n2624), .C(n2043), .D(n2495), .Y(n2622) );
  OAI22X1TS U2062 ( .A0(n2153), .A1(n10524), .B0(n2781), .B1(n2510), .Y(n2780)
         );
  OAI22X1TS U2036 ( .A0(n2057), .A1(n10592), .B0(n2073), .B1(n11525), .Y(n2745) );
  NOR2X1TS U2031 ( .A(n2740), .B(n2741), .Y(n1385) );
  INVX2TS U2029 ( .A(n1385), .Y(n1388) );
  OAI22X1TS U1884 ( .A0(n1672), .A1(n9765), .B0(n2012), .B1(n10954), .Y(n2570)
         );
  AOI22X1TS U1883 ( .A0(n10180), .A1(n11052), .B0(n11913), .B1(n12182), .Y(
        n2589) );
  AOI22X1TS U1870 ( .A0(n12186), .A1(n2577), .B0(n11051), .B1(n9749), .Y(n2573) );
  INVX2TS U1862 ( .A(n1465), .Y(n1466) );
  INVX2TS U1663 ( .A(n1360), .Y(n1359) );
  AOI22X1TS U1207 ( .A0(n1424), .A1(n1425), .B0(n1426), .B1(n1427), .Y(n1423)
         );
  OAI22X1TS U2203 ( .A0(n11147), .A1(n10208), .B0(n2095), .B1(n10280), .Y(
        n2921) );
  OAI22X1TS U2160 ( .A0(n12476), .A1(n10981), .B0(n11434), .B1(n9072), .Y(
        n2870) );
  INVX2TS U2147 ( .A(n1464), .Y(n1462) );
  OAI22X1TS U2128 ( .A0(n11126), .A1(n10216), .B0(n2121), .B1(n10256), .Y(
        n2845) );
  OAI22X1TS U2085 ( .A0(n12460), .A1(n10997), .B0(n11428), .B1(n9079), .Y(
        n2794) );
  OAI22X1TS U1185 ( .A0(n1389), .A1(n12756), .B0(n12692), .B1(n1390), .Y(N81)
         );
  AOI22X1TS U3550 ( .A0(n4023), .A1(n3354), .B0(n3355), .B1(n9126), .Y(n3933)
         );
  OAI22X1TS U3500 ( .A0(n3931), .A1(n12750), .B0(n12688), .B1(n3932), .Y(N228)
         );
  AOI22X1TS U1171 ( .A0(n12677), .A1(n1359), .B0(n1360), .B1(n9776), .Y(n1347)
         );
  AOI22X1TS U1820 ( .A0(n10184), .A1(n2514), .B0(n11537), .B1(n2494), .Y(n2458) );
  OAI211X1TS U1819 ( .A0(n1982), .A1(n2510), .B0(n2511), .C0(n2512), .Y(n2504)
         );
  OAI22X1TS U1818 ( .A0(n11555), .A1(n11531), .B0(n11459), .B1(n10593), .Y(
        n2505) );
  OAI22X1TS U1815 ( .A0(n10236), .A1(n12316), .B0(n11079), .B1(n11835), .Y(
        n2497) );
  AOI22X1TS U1799 ( .A0(n2469), .A1(n2058), .B0(n11561), .B1(n2470), .Y(n2467)
         );
  OAI211X1TS U1798 ( .A0(n2465), .A1(n2638), .B0(n2467), .C0(n2468), .Y(n2464)
         );
  OAI22X1TS U1165 ( .A0(n1345), .A1(n12755), .B0(n12692), .B1(n1346), .Y(N84)
         );
  AOI22X1TS U1849 ( .A0(n11500), .A1(n9087), .B0(n11955), .B1(n2549), .Y(n2547) );
  OAI211X1TS U1842 ( .A0(n2216), .A1(n10288), .B0(n2182), .C0(n2543), .Y(n2542) );
  AOI211X1TS U1841 ( .A0(n11823), .A1(n1682), .B0(n2541), .C0(n2542), .Y(n2515) );
  OAI22X1TS U1835 ( .A0(n10004), .A1(n10012), .B0(n9701), .B1(n11589), .Y(
        n2520) );
  OAI31X1TS U1826 ( .A0(n12359), .A1(n10584), .A2(n2518), .B0(n12180), .Y(
        n2517) );
  INVX2TS U1824 ( .A(n9242), .Y(n1382) );
  INVX2TS U1822 ( .A(n1455), .Y(n1454) );
  AOI22X1TS U1223 ( .A0(n9772), .A1(n1454), .B0(n1455), .B1(n9773), .Y(n1452)
         );
  AOI22X1TS U5433 ( .A0(n5823), .A1(n5148), .B0(n5149), .B1(n9318), .Y(n5730)
         );
  OAI22X1TS U5384 ( .A0(n5728), .A1(n12745), .B0(n12685), .B1(n5729), .Y(N164)
         );
  AOI22X1TS U5158 ( .A0(n5140), .A1(n5191), .B0(n5192), .B1(n9206), .Y(n5241)
         );
  OAI22X1TS U7014 ( .A0(n7002), .A1(n12738), .B0(n12691), .B1(n7003), .Y(N131)
         );
  AOI22X1TS U5982 ( .A0(n5823), .A1(n5231), .B0(n5232), .B1(n9317), .Y(n6323)
         );
  OAI22X1TS U5783 ( .A0(n6321), .A1(n12743), .B0(n12684), .B1(n6322), .Y(N161)
         );
  INVX2TS U2311 ( .A(n9083), .Y(n2229) );
  AOI22X1TS U2222 ( .A0(n2229), .A1(n1471), .B0(n1472), .B1(n9082), .Y(n2737)
         );
  OAI22X1TS U2024 ( .A0(n2735), .A1(n12753), .B0(n12690), .B1(n2736), .Y(N33)
         );
  AOI22X1TS U5062 ( .A0(n5131), .A1(n5132), .B0(n9203), .B1(n5133), .Y(n5129)
         );
  AOI22X1TS U1662 ( .A0(n2229), .A1(n1359), .B0(n1360), .B1(n9082), .Y(n2129)
         );
  OAI22X1TS U1611 ( .A0(n2127), .A1(n12753), .B0(n12691), .B1(n2128), .Y(N36)
         );
  OAI22X1TS U1147 ( .A0(n1306), .A1(n9039), .B0(n12693), .B1(n1307), .Y(N87)
         );
  AOI22X1TS U1295 ( .A0(n1465), .A1(n9270), .B0(n12672), .B1(n1466), .Y(n1523)
         );
  INVX2TS U1361 ( .A(n9239), .Y(n1386) );
  AOI22X1TS U1294 ( .A0(n1386), .A1(n9564), .B0(n9562), .B1(n9238), .Y(n1525)
         );
  OAI22X1TS U1289 ( .A0(n1521), .A1(n12754), .B0(n12691), .B1(n1522), .Y(N49)
         );
  AOI22X1TS U1266 ( .A0(n9269), .A1(n1448), .B0(n1449), .B1(n12672), .Y(n1500)
         );
  OAI22X1TS U1259 ( .A0(n1498), .A1(n12754), .B0(n12693), .B1(n1499), .Y(N51)
         );
  AOI22X1TS U1177 ( .A0(n1372), .A1(n9601), .B0(n9599), .B1(n9246), .Y(n1366)
         );
  OAI22X1TS U1172 ( .A0(n1362), .A1(n12755), .B0(n12693), .B1(n1363), .Y(N83)
         );
  AOI22X1TS U1229 ( .A0(n1465), .A1(n12666), .B0(n1437), .B1(n1466), .Y(n1459)
         );
  OAI22X1TS U1224 ( .A0(n1457), .A1(n12754), .B0(n12694), .B1(n1458), .Y(N65)
         );
  AOI22X1TS U1219 ( .A0(n12666), .A1(n1448), .B0(n1449), .B1(n1437), .Y(n1442)
         );
  OAI22X1TS U1214 ( .A0(n1440), .A1(n12756), .B0(n12693), .B1(n1441), .Y(N67)
         );
  AOI22X1TS U1163 ( .A0(n1338), .A1(n9611), .B0(n9609), .B1(n9254), .Y(n1337)
         );
  OAI22X1TS U1159 ( .A0(n1332), .A1(n12755), .B0(n12694), .B1(n1333), .Y(N85)
         );
  AOI22X1TS U1183 ( .A0(n1382), .A1(n9596), .B0(n9594), .B1(n9243), .Y(n1381)
         );
  OAI22X1TS U1179 ( .A0(n1376), .A1(n12756), .B0(n12692), .B1(n1377), .Y(N82)
         );
  AOI22X1TS U1464 ( .A0(n1774), .A1(n9426), .B0(n9427), .B1(n1776), .Y(N387)
         );
  AOI22X1TS U1387 ( .A0(n9140), .A1(n9319), .B0(n9320), .B1(n1628), .Y(N414)
         );
  AOI22X1TS U1382 ( .A0(n1619), .A1(n9412), .B0(n9413), .B1(n1621), .Y(N419)
         );
  AOI22X1TS U1390 ( .A0(n1633), .A1(n9327), .B0(n9328), .B1(n1635), .Y(N411)
         );
  AOI22X1TS U1381 ( .A0(n1616), .A1(n9408), .B0(n9409), .B1(n1618), .Y(N420)
         );
  AOI22X1TS U1389 ( .A0(n1630), .A1(n9323), .B0(n9324), .B1(n1632), .Y(N412)
         );
  AOI22X1TS U1343 ( .A0(n9174), .A1(n9389), .B0(n9390), .B1(n9173), .Y(N454)
         );
  AOI22X1TS U1351 ( .A0(n9168), .A1(n9304), .B0(n9305), .B1(n9167), .Y(N446)
         );
  AOI22X1TS U1405 ( .A0(n9274), .A1(n9614), .B0(n9615), .B1(n9273), .Y(N401)
         );
  AOI22X1TS U1395 ( .A0(n1385), .A1(n9590), .B0(n9591), .B1(n1388), .Y(N406)
         );
  AOI22X1TS U1269 ( .A0(n1396), .A1(n9548), .B0(n9549), .B1(n1397), .Y(N502)
         );
  AOI22X1TS U1359 ( .A0(n1386), .A1(n9577), .B0(n9578), .B1(n9238), .Y(N438)
         );
  AOI22X1TS U1471 ( .A0(n1785), .A1(n9336), .B0(n9337), .B1(n1787), .Y(N380)
         );
  AOI22X1TS U1399 ( .A0(n1352), .A1(n9599), .B0(n9600), .B1(n1353), .Y(N404)
         );
  AOI22X1TS U1282 ( .A0(n1512), .A1(n9464), .B0(n9465), .B1(n1513), .Y(N494)
         );
  AOI22X1TS U1335 ( .A0(n1558), .A1(n9478), .B0(n9479), .B1(n1560), .Y(N462)
         );
  AOI22X1TS U1371 ( .A0(n1598), .A1(n9493), .B0(n9494), .B1(n1600), .Y(N430)
         );
  AOI211X1TS U7799 ( .A0(n12625), .A1(n8197), .B0(n8198), .C0(n8199), .Y(n8196) );
  AOI211X1TS U7721 ( .A0(n12108), .A1(n11886), .B0(n7941), .C0(n8130), .Y(
        n8128) );
  NOR2X1TS U7716 ( .A(n11939), .B(n12108), .Y(n7927) );
  AOI211X1TS U7607 ( .A0(n11854), .A1(n12371), .B0(n7687), .C0(n8035), .Y(
        n8033) );
  OAI22X1TS U7229 ( .A0(n1513), .A1(n1296), .B0(n9784), .B1(n1512), .Y(n7018)
         );
  OAI22X1TS U7152 ( .A0(n7123), .A1(n12465), .B0(n7263), .B1(n12122), .Y(n7262) );
  OAI22X1TS U7274 ( .A0(n10034), .A1(n12465), .B0(n10677), .B1(n10054), .Y(
        n7538) );
  AOI22X1TS U1136 ( .A0(n1284), .A1(n1285), .B0(n1286), .B1(n1287), .Y(n1283)
         );
  AOI22X1TS U7528 ( .A0(n11886), .A1(n11940), .B0(n11812), .B1(n12108), .Y(
        n7938) );
  AOI211X1TS U7411 ( .A0(n11546), .A1(n10669), .B0(n7796), .C0(n7053), .Y(
        n7795) );
  AOI211X1TS U8705 ( .A0(n12108), .A1(n11048), .B0(n8662), .C0(n8663), .Y(
        n8661) );
  AOI211X1TS U4059 ( .A0(n11224), .A1(n10773), .B0(n4689), .C0(n4690), .Y(
        n4688) );
  AOI211X1TS U4057 ( .A0(n11985), .A1(n11285), .B0(n4685), .C0(n4686), .Y(
        n4684) );
  AOI211X1TS U4079 ( .A0(n11988), .A1(n12580), .B0(n4708), .C0(n4709), .Y(
        n4706) );
  AOI211X1TS U3984 ( .A0(n11230), .A1(n10761), .B0(n4617), .C0(n4618), .Y(
        n4616) );
  AOI211X1TS U3982 ( .A0(n12000), .A1(n11332), .B0(n4613), .C0(n4614), .Y(
        n4612) );
  NOR2X1TS U4265 ( .A(n12490), .B(n12208), .Y(n4867) );
  AOI211X1TS U4224 ( .A0(n10395), .A1(n12029), .B0(n4832), .C0(n4498), .Y(
        n4831) );
  NOR2X1TS U4357 ( .A(n12377), .B(n10159), .Y(n4758) );
  AOI31X1TS U4352 ( .A0(n10163), .A1(n12039), .A2(n9664), .B0(n12065), .Y(
        n4918) );
  NOR2X1TS U4330 ( .A(n11798), .B(n11786), .Y(n4276) );
  AOI31X1TS U4327 ( .A0(n3517), .A1(n10945), .A2(n12065), .B0(n11803), .Y(
        n4901) );
  AOI211X1TS U4324 ( .A0(n11273), .A1(n4900), .B0(n4901), .C0(n4371), .Y(n4899) );
  AOI211X1TS U3362 ( .A0(n4131), .A1(n10476), .B0(n3587), .C0(n3588), .Y(n3585) );
  AOI211X1TS U5942 ( .A0(n11413), .A1(n11007), .B0(n6489), .C0(n6490), .Y(
        n6488) );
  AOI211X1TS U5940 ( .A0(n12047), .A1(n11317), .B0(n6485), .C0(n6486), .Y(
        n6484) );
  AOI211X1TS U5867 ( .A0(n11407), .A1(n10995), .B0(n6417), .C0(n6418), .Y(
        n6416) );
  AOI211X1TS U5865 ( .A0(n12033), .A1(n11269), .B0(n6413), .C0(n6414), .Y(
        n6412) );
  AOI211X1TS U5887 ( .A0(n12036), .A1(n12583), .B0(n6436), .C0(n6437), .Y(
        n6434) );
  OAI32X1TS U6140 ( .A0(n10940), .A1(n6662), .A2(n12055), .B0(n12281), .B1(
        n6662), .Y(n6660) );
  NOR2X1TS U6118 ( .A(n11349), .B(n12278), .Y(n6311) );
  AOI211X1TS U6111 ( .A0(n11723), .A1(n9407), .B0(n6636), .C0(n6365), .Y(n6635) );
  NOR2X1TS U6239 ( .A(n12449), .B(n10141), .Y(n6558) );
  AOI31X1TS U6234 ( .A0(n10412), .A1(n11978), .A2(n9762), .B0(n12198), .Y(
        n6717) );
  NOR2X1TS U6212 ( .A(n11684), .B(n11675), .Y(n6043) );
  AOI211X1TS U7450 ( .A0(n11615), .A1(n12371), .B0(n7857), .C0(n7858), .Y(
        n7856) );
  AOI211X1TS U3385 ( .A0(n12031), .A1(n10877), .B0(n3645), .C0(n3646), .Y(
        n3642) );
  AOI211X1TS U6408 ( .A0(n11276), .A1(n9364), .B0(n6770), .C0(n6771), .Y(n6769) );
  AOI211X1TS U6781 ( .A0(n11724), .A1(n12294), .B0(n6886), .C0(n6887), .Y(
        n6885) );
  AOI211X1TS U6044 ( .A0(n11696), .A1(n10951), .B0(n6578), .C0(n6579), .Y(
        n6576) );
  AOI211X1TS U4525 ( .A0(n11327), .A1(n9157), .B0(n4971), .C0(n4972), .Y(n4970) );
  AOI211X1TS U4161 ( .A0(n12073), .A1(n10799), .B0(n4778), .C0(n4779), .Y(
        n4776) );
  AOI22X1TS U7444 ( .A0(n9865), .A1(n11517), .B0(n11617), .B1(n12617), .Y(
        n7844) );
  AOI211X1TS U7429 ( .A0(n12616), .A1(n10729), .B0(n7816), .C0(n7633), .Y(
        n7814) );
  AOI22X1TS U6954 ( .A0(n6941), .A1(n1641), .B0(n1643), .B1(n6942), .Y(n6940)
         );
  NOR2X1TS U7370 ( .A(n11598), .B(n11868), .Y(n7741) );
  AOI22X1TS U7050 ( .A0(n6935), .A1(n7028), .B0(n9212), .B1(n1528), .Y(n7026)
         );
  AOI211X1TS U6603 ( .A0(n11324), .A1(n9371), .B0(n6828), .C0(n6829), .Y(n6827) );
  AOI211X1TS U4720 ( .A0(n11279), .A1(n9166), .B0(n5029), .C0(n5030), .Y(n5028) );
  OAI22X1TS U4028 ( .A0(n9655), .A1(n12428), .B0(n9162), .B1(n11292), .Y(n4655) );
  OAI22X1TS U3953 ( .A0(n9658), .A1(n12444), .B0(n9153), .B1(n11340), .Y(n4583) );
  AOI211X1TS U3836 ( .A0(n11988), .A1(n11225), .B0(n4136), .C0(n4435), .Y(
        n4434) );
  AOI22X1TS U3896 ( .A0(n10391), .A1(n10808), .B0(n12199), .B1(n11214), .Y(
        n4511) );
  OAI22X1TS U3266 ( .A0(n1596), .A1(n9131), .B0(n3330), .B1(n9092), .Y(n3408)
         );
  AOI211X1TS U3800 ( .A0(n12000), .A1(n11231), .B0(n4080), .C0(n4395), .Y(
        n4394) );
  OAI22X1TS U5148 ( .A0(n1582), .A1(n9143), .B0(n5124), .B1(n9279), .Y(n5205)
         );
  NOR2X1TS U2960 ( .A(n9627), .B(n10240), .Y(n2297) );
  NOR2X1TS U2763 ( .A(n12599), .B(n10263), .Y(n2364) );
  AOI22X1TS U2729 ( .A0(n11136), .A1(n10538), .B0(n12137), .B1(n12598), .Y(
        n3196) );
  AOI31X1TS U2454 ( .A0(n9927), .A1(n12563), .A2(n9960), .B0(n12159), .Y(n3116) );
  NOR2X1TS U2446 ( .A(n12359), .B(n12192), .Y(n3089) );
  OAI22X1TS U1893 ( .A0(n9999), .A1(n12562), .B0(n10602), .B1(n9964), .Y(n2602) );
  AOI211X1TS U1538 ( .A0(n12110), .A1(n1961), .B0(n1962), .C0(n1963), .Y(n1958) );
  NOR2X1TS U1533 ( .A(n9972), .B(n12133), .Y(n1757) );
  NOR2X1TS U1509 ( .A(n9984), .B(n12147), .Y(n1719) );
  AOI211X1TS U2171 ( .A0(n10272), .A1(n11846), .B0(n2411), .C0(n2894), .Y(
        n2893) );
  NOR2X1TS U2427 ( .A(n11822), .B(n11912), .Y(n2552) );
  AOI211X1TS U1852 ( .A0(n12325), .A1(n10679), .B0(n2555), .C0(n2556), .Y(
        n2554) );
  AOI211X1TS U5823 ( .A0(n11331), .A1(n12299), .B0(n6376), .C0(n6377), .Y(
        n6375) );
  AOI211X1TS U3676 ( .A0(n11732), .A1(n12580), .B0(n3754), .C0(n4227), .Y(
        n4226) );
  AOI22X1TS U5778 ( .A0(n12055), .A1(n12279), .B0(n12062), .B1(n11742), .Y(
        n6313) );
  AOI211X1TS U5776 ( .A0(n11741), .A1(n10177), .B0(n6309), .C0(n6310), .Y(
        n6308) );
  AOI211X1TS U5771 ( .A0(n11742), .A1(n10947), .B0(n5570), .C0(n6305), .Y(
        n6304) );
  AOI211X1TS U5718 ( .A0(n12047), .A1(n11414), .B0(n5936), .C0(n6238), .Y(
        n6237) );
  AOI211X1TS U7170 ( .A0(n11856), .A1(n12141), .B0(n7323), .C0(n7324), .Y(
        n7320) );
  AOI211X1TS U1710 ( .A0(n12296), .A1(n12600), .B0(n2325), .C0(n2326), .Y(
        n2320) );
  OAI22X1TS U5911 ( .A0(n9719), .A1(n12399), .B0(n9368), .B1(n11313), .Y(n6455) );
  AOI211X1TS U5682 ( .A0(n12033), .A1(n11408), .B0(n5880), .C0(n6198), .Y(
        n6197) );
  OAI22X1TS U2345 ( .A0(n10523), .A1(n11858), .B0(n10631), .B1(n10626), .Y(
        n3037) );
  AOI211X1TS U1675 ( .A0(n12302), .A1(n12604), .B0(n2258), .C0(n2259), .Y(
        n2253) );
  OAI22X1TS U2521 ( .A0(n10955), .A1(n12562), .B0(n10684), .B1(n9700), .Y(
        n3132) );
  AOI22X1TS U1239 ( .A0(n1480), .A1(n1417), .B0(n1420), .B1(n9227), .Y(n1479)
         );
  OAI22X1TS U2889 ( .A0(n2725), .A1(n12461), .B0(n2272), .B1(n10575), .Y(n3247) );
  AOI211X1TS U2869 ( .A0(n10579), .A1(n12367), .B0(n1748), .C0(n3243), .Y(
        n3242) );
  OAI22X1TS U2817 ( .A0(n2423), .A1(n12458), .B0(n2279), .B1(n11470), .Y(n3219) );
  NOR2X1TS U2814 ( .A(n10565), .B(n12367), .Y(n2244) );
  AOI221X1TS U2291 ( .A0(n12187), .A1(n2222), .B0(n12194), .B1(n2201), .C0(
        n2999), .Y(n2968) );
  AOI211X1TS U2253 ( .A0(n12154), .A1(n2185), .B0(n2186), .C0(n2965), .Y(n2964) );
  OAI22X1TS U2692 ( .A0(n2692), .A1(n12474), .B0(n2339), .B1(n10548), .Y(n3187) );
  AOI211X1TS U2672 ( .A0(n10551), .A1(n12374), .B0(n1710), .C0(n3183), .Y(
        n3182) );
  AOI22X1TS U1410 ( .A0(n9784), .A1(n9507), .B0(n9508), .B1(n1296), .Y(N398)
         );
  AOI22X1TS U3189 ( .A0(n3346), .A1(n1633), .B0(n1635), .B1(n9188), .Y(n3343)
         );
  AOI22X1TS U5067 ( .A0(n5140), .A1(n1619), .B0(n1621), .B1(n9207), .Y(n5136)
         );
  AOI22X1TS U3210 ( .A0(n3372), .A1(n9140), .B0(n1628), .B1(n1549), .Y(n3369)
         );
  AOI22X1TS U5088 ( .A0(n5166), .A1(n1612), .B0(n1614), .B1(n1534), .Y(n5163)
         );
  AOI22X1TS U2003 ( .A0(n10240), .A1(n10561), .B0(n12130), .B1(n9057), .Y(
        n2721) );
  AOI22X1TS U1961 ( .A0(n10264), .A1(n10533), .B0(n12144), .B1(n9064), .Y(
        n2688) );
  AOI211X1TS U1910 ( .A0(n11560), .A1(n12308), .B0(n2146), .C0(n2627), .Y(
        n2626) );
  AOI22X1TS U1152 ( .A0(n1315), .A1(n9270), .B0(n12672), .B1(n9265), .Y(n1308)
         );
  AOI22X1TS U1263 ( .A0(n9772), .A1(n1382), .B0(n9242), .B1(n1456), .Y(n1503)
         );
  AOI32XLTS U1119 ( .A0(dcnt[1]), .A1(n1262), .A2(dcnt[0]), .B0(n1263), .B1(
        n1262), .Y(n1261) );
  NOR4XLTS U7208 ( .A(n7409), .B(n7410), .C(n7411), .D(n7412), .Y(n7151) );
  NOR4XLTS U8450 ( .A(n7865), .B(n7118), .C(n8563), .D(n8564), .Y(n7346) );
  AOI22X1TS U7875 ( .A0(n11862), .A1(n11591), .B0(n11125), .B1(n11145), .Y(
        n8282) );
  NOR4XLTS U8635 ( .A(n7911), .B(n8629), .C(n8630), .D(n8631), .Y(n7198) );
  NOR4XLTS U3432 ( .A(n3777), .B(n3778), .C(n3779), .D(n3780), .Y(n3564) );
  NOR4XLTS U3407 ( .A(n3711), .B(n3712), .C(n3713), .D(n3714), .Y(n3525) );
  AOI22X1TS U4329 ( .A0(n10155), .A1(n11786), .B0(n11792), .B1(n10800), .Y(
        n4898) );
  NOR4XLTS U5303 ( .A(n5532), .B(n5533), .C(n5534), .D(n5535), .Y(n5362) );
  NOR4XLTS U5278 ( .A(n5466), .B(n5467), .C(n5468), .D(n5469), .Y(n5323) );
  AOI22X1TS U7227 ( .A0(n6926), .A1(n1282), .B0(n7018), .B1(n9794), .Y(n7342)
         );
  NOR4XLTS U5338 ( .A(n5618), .B(n5619), .C(n5620), .D(n5621), .Y(n5277) );
  NOR4XLTS U6753 ( .A(n6864), .B(n6865), .C(n6866), .D(n6867), .Y(n5644) );
  NOR4XLTS U7442 ( .A(n7839), .B(n7840), .C(n7841), .D(n7842), .Y(n7305) );
  OAI32X1TS U7554 ( .A0(n7973), .A1(n11171), .A2(n12642), .B0(n12470), .B1(
        n7973), .Y(n7971) );
  NOR4XLTS U3456 ( .A(n3823), .B(n3824), .C(n3825), .D(n3826), .Y(n3479) );
  AOI22X1TS U3863 ( .A0(n12238), .A1(n12053), .B0(n11279), .B1(n10778), .Y(
        n4463) );
  NOR4XLTS U3853 ( .A(n4446), .B(n4447), .C(n4448), .D(n4449), .Y(n3878) );
  AOI22X1TS U2926 ( .A0(n11116), .A1(n10564), .B0(n12123), .B1(n12602), .Y(
        n3256) );
  NOR4XLTS U1885 ( .A(n2591), .B(n2592), .C(n2593), .D(n2594), .Y(n2006) );
  NOR4XLTS U2038 ( .A(n2751), .B(n2752), .C(n1953), .D(n2753), .Y(n2132) );
  OAI32X1TS U2066 ( .A0(n10962), .A1(n9681), .A2(n9951), .B0(n11460), .B1(
        n10961), .Y(n2789) );
  NOR4XLTS U2063 ( .A(n2782), .B(n2783), .C(n2784), .D(n2785), .Y(n1952) );
  NOR4XLTS U2359 ( .A(n2137), .B(n2751), .C(n3052), .D(n3053), .Y(n1959) );
  AOI22X1TS U1722 ( .A0(n9744), .A1(n10971), .B0(n10271), .B1(n10299), .Y(
        n2343) );
  NOR4XLTS U5735 ( .A(n6249), .B(n6250), .C(n6251), .D(n6252), .Y(n5708) );
  AOI22X1TS U3260 ( .A0(n3428), .A1(n12665), .B0(n3408), .B1(n3429), .Y(n3425)
         );
  AOI22X1TS U3258 ( .A0(n9168), .A1(n9321), .B0(n9319), .B1(n9167), .Y(n3427)
         );
  AOI22X1TS U5140 ( .A0(n9174), .A1(n9406), .B0(n9404), .B1(n9173), .Y(n5224)
         );
  AOI22X1TS U3249 ( .A0(n12665), .A1(n3415), .B0(n3416), .B1(n3408), .Y(n3412)
         );
  AOI22X1TS U5130 ( .A0(n12664), .A1(n5212), .B0(n5213), .B1(n5205), .Y(n5209)
         );
  AOI22X1TS U6983 ( .A0(n1305), .A1(n6972), .B0(n1597), .B1(n9780), .Y(n6971)
         );
  NOR4XLTS U2339 ( .A(n3036), .B(n3037), .C(n3038), .D(n3039), .Y(n2743) );
  AOI22X1TS U2135 ( .A0(n12126), .A1(n12130), .B0(n10560), .B1(n10988), .Y(
        n2851) );
  NOR4XLTS U2497 ( .A(n3131), .B(n3132), .C(n3133), .D(n3134), .Y(n2588) );
  AOI22X1TS U2210 ( .A0(n12137), .A1(n12145), .B0(n10532), .B1(n10971), .Y(
        n2927) );
  AOI22X1TS U6995 ( .A0(n6980), .A1(n6926), .B0(n9793), .B1(n9127), .Y(n6979)
         );
  AOI22X1TS U1151 ( .A0(n9274), .A1(n9621), .B0(n9619), .B1(n9273), .Y(n1311)
         );
  NOR4XLTS U7834 ( .A(n8241), .B(n8242), .C(n8243), .D(n8244), .Y(n7468) );
  INVX2TS U7231 ( .A(n9783), .Y(n1296) );
  NOR3X1TS U8474 ( .A(sa13[6]), .B(n8578), .C(n12084), .Y(n7510) );
  AOI32X1TS U5228 ( .A0(sa12[0]), .A1(n10852), .A2(n5327), .B0(n10421), .B1(
        n10853), .Y(n5325) );
  AOI22X1TS U1141 ( .A0(n9784), .A1(n9466), .B0(n9464), .B1(n1296), .Y(n1293)
         );
  INVX2TS U3313 ( .A(n9140), .Y(n1628) );
  INVX2TS U3297 ( .A(n9137), .Y(n1632) );
  INVX2TS U5178 ( .A(n9149), .Y(n1618) );
  INVX2TS U3216 ( .A(n9085), .Y(n1625) );
  INVX2TS U5096 ( .A(n9272), .Y(n1611) );
  NOR4XLTS U8280 ( .A(n8226), .B(n7442), .C(n8511), .D(n8512), .Y(n7957) );
  NOR4XLTS U5507 ( .A(n5648), .B(n5942), .C(n5943), .D(n5944), .Y(n1771) );
  NOR4XLTS U5361 ( .A(n5678), .B(n5679), .C(n5680), .D(n5681), .Y(n5247) );
  NOR4XLTS U1701 ( .A(n1848), .B(n2298), .C(n2299), .D(n2300), .Y(n1433) );
  NOR4XLTS U4887 ( .A(n5076), .B(n4317), .C(n5077), .D(n5078), .Y(n4468) );
  NOR4XLTS U1513 ( .A(n1889), .B(n1890), .C(n1891), .D(n1892), .Y(n1486) );
  NOR4XLTS U7697 ( .A(n7043), .B(n7156), .C(n8102), .D(n8103), .Y(n6990) );
  NOR4XLTS U7397 ( .A(n7773), .B(n7774), .C(n7775), .D(n7776), .Y(n7023) );
  NOR4XLTS U5373 ( .A(n5703), .B(n5704), .C(n5705), .D(n5706), .Y(n5196) );
  NOR4XLTS U2784 ( .A(n2705), .B(n2446), .C(n3202), .D(n3203), .Y(n1395) );
  NOR4XLTS U2980 ( .A(n2624), .B(n2476), .C(n2063), .D(n3262), .Y(n1399) );
  NOR4XLTS U6742 ( .A(n5989), .B(n6856), .C(n6857), .D(n6858), .Y(n5174) );
  NOR4XLTS U3490 ( .A(n3898), .B(n3899), .C(n3900), .D(n3901), .Y(n3337) );
  NOR4XLTS U5750 ( .A(n5979), .B(n5951), .C(n6270), .D(n6271), .Y(n5157) );
  NOR4XLTS U4859 ( .A(n5057), .B(n5058), .C(n5059), .D(n5060), .Y(n3379) );
  NOR4XLTS U3868 ( .A(n4287), .B(n3898), .C(n4328), .D(n4467), .Y(n3363) );
  CLKBUFX2TS U8228 ( .A(sa31[5]), .Y(n8453) );
  CLKBUFX2TS U8216 ( .A(sa31[2]), .Y(n7656) );
  CLKINVX2TS U6940 ( .A(sa01[5]), .Y(n6918) );
  CLKINVX2TS U8225 ( .A(sa31[0]), .Y(n8467) );
  INVX1TS U1880 ( .A(sa32[1]), .Y(n2558) );
  INVX2TS U5045 ( .A(sa00[1]), .Y(n4515) );
  CLKINVX2TS U8414 ( .A(sa02[5]), .Y(n8546) );
  NOR2X1TS U1122 ( .A(dcnt[0]), .B(dcnt[1]), .Y(n1263) );
  INVX2TS U8608 ( .A(sa13[1]), .Y(n7528) );
  CLKBUFX2TS U2951 ( .A(sa10[0]), .Y(n1769) );
  INVX2TS U2975 ( .A(sa10[6]), .Y(n2430) );
  INVX2TS U2972 ( .A(sa10[2]), .Y(n2274) );
  INVX2TS U2778 ( .A(sa21[6]), .Y(n2386) );
  CLKBUFX2TS U8400 ( .A(sa02[4]), .Y(n7991) );
  CLKBUFX2TS U2754 ( .A(sa21[0]), .Y(n1731) );
  INVX2TS U2775 ( .A(sa21[2]), .Y(n2341) );
  CLKINVX1TS U1121 ( .A(n1260), .Y(n1264) );
  NAND3XLTS U5090 ( .A(n133), .B(n139), .C(n12667), .Y(n5167) );
  NOR2X1TS U2552 ( .A(sa32[0]), .B(n10354), .Y(n2996) );
  INVX2TS U2583 ( .A(n10088), .Y(n2997) );
  INVX2TS U5040 ( .A(n9788), .Y(n5112) );
  NOR2X1TS U4838 ( .A(sa22[1]), .B(n10084), .Y(n5052) );
  AND2X2TS U2555 ( .A(n10088), .B(sa32[5]), .Y(n2029) );
  NOR2X1TS U4841 ( .A(n9447), .B(n9840), .Y(n5034) );
  INVX2TS U6348 ( .A(n9812), .Y(n6049) );
  NOR2X1TS U4853 ( .A(n11190), .B(n9451), .Y(n4697) );
  NOR2X1TS U2959 ( .A(sa10[2]), .B(n10699), .Y(n2838) );
  INVX2TS U4465 ( .A(n9888), .Y(n4282) );
  NOR2X1TS U6281 ( .A(n9808), .B(n10709), .Y(n6719) );
  NOR2X1TS U5037 ( .A(n10314), .B(sa00[1]), .Y(n5106) );
  INVX2TS U3158 ( .A(n10096), .Y(n2652) );
  NOR2X1TS U2562 ( .A(sa32[7]), .B(n9848), .Y(n3138) );
  AND2X2TS U4848 ( .A(n11191), .B(n9451), .Y(n4197) );
  INVX2TS U3143 ( .A(n9530), .Y(n3306) );
  NOR2X1TS U2520 ( .A(n9852), .B(sa32[1]), .Y(n3130) );
  OR2X2TS U8413 ( .A(n8546), .B(n9832), .Y(n8237) );
  OR2X2TS U3135 ( .A(n9522), .B(n9856), .Y(n3305) );
  NOR2X1TS U4828 ( .A(n9458), .B(sa22[5]), .Y(n5033) );
  NOR2X1TS U8421 ( .A(sa02[2]), .B(sa02[4]), .Y(n8525) );
  INVX2TS U2578 ( .A(n10349), .Y(n2035) );
  AND2X2TS U4835 ( .A(sa22[1]), .B(n10084), .Y(n4692) );
  NOR2X1TS U6306 ( .A(sa30[6]), .B(n9812), .Y(n6724) );
  AND2X2TS U4440 ( .A(n10748), .B(n9888), .Y(n4281) );
  INVX2TS U2950 ( .A(n10028), .Y(n2113) );
  INVX2TS U4857 ( .A(n9458), .Y(n3568) );
  INVX2TS U3147 ( .A(n9522), .Y(n2660) );
  INVX2TS U2577 ( .A(sa32[4]), .Y(n3139) );
  NOR2X1TS U3155 ( .A(n10359), .B(n10364), .Y(n3322) );
  INVX2TS U2584 ( .A(n10355), .Y(n2599) );
  NOR2X1TS U3129 ( .A(sa03[2]), .B(sa03[4]), .Y(n3313) );
  OR2X2TS U5051 ( .A(n10318), .B(n5116), .Y(n4570) );
  AND2X2TS U5031 ( .A(n10313), .B(n4515), .Y(n4545) );
  OR2X2TS U2558 ( .A(n10350), .B(n9844), .Y(n3100) );
  INVX2TS U4847 ( .A(n10080), .Y(n4464) );
  INVX2TS U2575 ( .A(n9852), .Y(n3002) );
  AND2X2TS U6351 ( .A(n10715), .B(n9820), .Y(n6565) );
  NOR2X1TS U4400 ( .A(n9884), .B(n10742), .Y(n4920) );
  AND2X2TS U2955 ( .A(n2430), .B(n9282), .Y(n2454) );
  AND2X2TS U8578 ( .A(n11196), .B(n7528), .Y(n7546) );
  AND2X2TS U2758 ( .A(n2386), .B(sa21[1]), .Y(n2410) );
  NOR2X1TS U8556 ( .A(n9860), .B(n10738), .Y(n8611) );
  AND2X2TS U8589 ( .A(n9876), .B(n9872), .Y(n8050) );
  OR2X2TS U8560 ( .A(n9868), .B(n9864), .Y(n7905) );
  NOR2X1TS U4643 ( .A(sa11[1]), .B(n10056), .Y(n4994) );
  AND2X2TS U4640 ( .A(sa11[1]), .B(n10056), .Y(n4620) );
  INVX2TS U6740 ( .A(n9545), .Y(n5366) );
  NOR2X1TS U4658 ( .A(n11168), .B(sa11[4]), .Y(n4625) );
  AND2X2TS U6523 ( .A(sa12[1]), .B(n10076), .Y(n6420) );
  NOR2X1TS U8186 ( .A(n9366), .B(n10340), .Y(n8470) );
  INVX2TS U4662 ( .A(n9358), .Y(n3529) );
  NOR2X1TS U6736 ( .A(n11201), .B(n9538), .Y(n6497) );
  INVX2TS U8204 ( .A(n10336), .Y(n7730) );
  OR2X2TS U8605 ( .A(sa13[1]), .B(n11197), .Y(n8580) );
  NOR2X1TS U6721 ( .A(sa23[1]), .B(n10104), .Y(n6851) );
  NOR2X1TS U8394 ( .A(sa02[7]), .B(sa02[5]), .Y(n8535) );
  INVX2TS U6730 ( .A(n10100), .Y(n6267) );
  NOR2X1TS U4425 ( .A(n10747), .B(n9888), .Y(n4925) );
  AND2X2TS U8774 ( .A(n9804), .B(n9800), .Y(n8116) );
  NOR2X1TS U8368 ( .A(n10732), .B(n11174), .Y(n8539) );
  NOR2X1TS U6902 ( .A(sa01[0]), .B(sa01[3]), .Y(n6910) );
  OR2X2TS U6937 ( .A(n6917), .B(n10048), .Y(n6302) );
  INVX2TS U6923 ( .A(n9824), .Y(n6318) );
  AND2X2TS U4653 ( .A(n11168), .B(n9351), .Y(n4153) );
  NOR2X1TS U6526 ( .A(sa12[1]), .B(n10076), .Y(n6793) );
  INVX2TS U2753 ( .A(n10060), .Y(n2087) );
  NOR2X1TS U8383 ( .A(n10345), .B(n11181), .Y(n8520) );
  AND2X2TS U6731 ( .A(n11201), .B(n9538), .Y(n6107) );
  INVX2TS U6535 ( .A(n10072), .Y(n6227) );
  NOR2X1TS U6541 ( .A(n11185), .B(n9435), .Y(n6425) );
  NOR2X1TS U6921 ( .A(n10722), .B(sa01[5]), .Y(n6891) );
  AND2X2TS U6718 ( .A(sa23[1]), .B(n10104), .Y(n6492) );
  OR2X2TS U8746 ( .A(n9796), .B(sa20[2]), .Y(n7952) );
  NOR2X1TS U6529 ( .A(sa12[3]), .B(sa12[0]), .Y(n6775) );
  AND2X2TS U6536 ( .A(n11186), .B(n9435), .Y(n6063) );
  NOR2X1TS U6891 ( .A(sa01[6]), .B(n9824), .Y(n6906) );
  NOR2X1TS U6711 ( .A(n9545), .B(n9541), .Y(n6832) );
  NOR2X1TS U6516 ( .A(sa12[7]), .B(n9439), .Y(n6774) );
  INVX2TS U6545 ( .A(sa12[7]), .Y(n5327) );
  NOR2X1TS U8742 ( .A(n9792), .B(n10704), .Y(n8676) );
  INVX2TS U4652 ( .A(n10052), .Y(n4424) );
  NOR2X1TS U4646 ( .A(n9348), .B(n9828), .Y(n4976) );
  AND2X2TS U4468 ( .A(n10752), .B(n9896), .Y(n4765) );
  OR2X2TS U8791 ( .A(n9286), .B(sa20[6]), .Y(n8649) );
  INVX2TS U8795 ( .A(n10040), .Y(n8644) );
  INVX2TS U8401 ( .A(n10068), .Y(n8540) );
  OR2X2TS U8181 ( .A(n10335), .B(sa31[2]), .Y(n8341) );
  NOR2X1TS U2762 ( .A(sa21[2]), .B(n10726), .Y(n2914) );
  NOR2X1TS U6724 ( .A(n9534), .B(sa23[0]), .Y(n6833) );
  INVX2TS U8749 ( .A(n9286), .Y(n7440) );
  NOR2X1TS U4633 ( .A(n9358), .B(n9355), .Y(n4975) );
  OR4X2TS U8536 ( .A(sa13[0]), .B(n10738), .C(sa13[7]), .D(sa13[5]), .Y(n7106)
         );
  OR2X2TS U8399 ( .A(n8540), .B(n9881), .Y(n7988) );
  AND3X2TS U8307 ( .A(n10731), .B(n11174), .C(n8525), .Y(n7446) );
  CLKINVX2TS U8223 ( .A(n8463), .Y(n8454) );
  CLKAND2X2TS U2865 ( .A(n2864), .B(n3241), .Y(n1939) );
  NOR3X1TS U8391 ( .A(n10732), .B(sa02[1]), .C(n9882), .Y(n8180) );
  OR2X2TS U4856 ( .A(n3568), .B(n9454), .Y(n4439) );
  OR2X2TS U8371 ( .A(sa02[4]), .B(n8540), .Y(n7619) );
  INVX1TS U6530 ( .A(n5693), .Y(n6797) );
  OR2X2TS U3146 ( .A(n2660), .B(n9855), .Y(n3075) );
  CLKINVX1TS U3113 ( .A(n3313), .Y(n2661) );
  AND2X2TS U6534 ( .A(n6227), .B(n10076), .Y(n6747) );
  AND2X2TS U6513 ( .A(n9439), .B(n5327), .Y(n5830) );
  AND2X2TS U4651 ( .A(n4424), .B(n10056), .Y(n4948) );
  CLKINVX2TS U6735 ( .A(n6497), .Y(n6268) );
  NOR2XLTS U6117 ( .A(n10048), .B(n6640), .Y(n5677) );
  OR2X2TS U5022 ( .A(n5112), .B(n9278), .Y(n5102) );
  INVX1TS U6725 ( .A(n5718), .Y(n6855) );
  NOR2XLTS U8236 ( .A(n11181), .B(n8488), .Y(n8211) );
  AND2X2TS U4630 ( .A(n9355), .B(n3529), .Y(n4030) );
  AND2X2TS U6708 ( .A(n9541), .B(n5366), .Y(n5886) );
  INVX1TS U4647 ( .A(n3863), .Y(n4998) );
  CLKINVX2TS U4657 ( .A(n4625), .Y(n4425) );
  OR2X2TS U6739 ( .A(n5366), .B(sa23[5]), .Y(n6242) );
  OR2X2TS U8205 ( .A(n10340), .B(n9365), .Y(n8452) );
  OR2X2TS U8202 ( .A(n7730), .B(n9854), .Y(n7727) );
  CLKINVX1TS U5043 ( .A(n5103), .Y(n5115) );
  AND2X2TS U3112 ( .A(n9856), .B(n2660), .Y(n2163) );
  OR2X2TS U4661 ( .A(n3529), .B(sa11[5]), .Y(n4399) );
  OR2X2TS U6544 ( .A(n5327), .B(sa12[5]), .Y(n6202) );
  NAND2XLTS U2288 ( .A(n2996), .B(n2997), .Y(n2617) );
  OR2X2TS U8187 ( .A(n10335), .B(n9853), .Y(n7694) );
  AND2X2TS U3173 ( .A(n10360), .B(n10363), .Y(n2651) );
  AND2X2TS U3122 ( .A(n3306), .B(sa03[7]), .Y(n2748) );
  CLKINVX2TS U6540 ( .A(n6425), .Y(n6228) );
  AND2X2TS U6729 ( .A(n6267), .B(n10104), .Y(n6805) );
  INVX1TS U4974 ( .A(n4516), .Y(n4876) );
  AND2X2TS U8794 ( .A(n8644), .B(n9286), .Y(n8641) );
  INVX1TS U2978 ( .A(n3249), .Y(n2112) );
  NOR2XLTS U5379 ( .A(n9534), .B(n5718), .Y(n5392) );
  INVX1TS U2781 ( .A(n3189), .Y(n2086) );
  AND2X2TS U2973 ( .A(n2430), .B(n9281), .Y(n2822) );
  AND2X2TS U4451 ( .A(n10753), .B(n9895), .Y(n4246) );
  CLKINVX2TS U2761 ( .A(n2914), .Y(n3185) );
  INVX1TS U4842 ( .A(n3888), .Y(n5056) );
  CLKINVX2TS U4852 ( .A(n4697), .Y(n4465) );
  OR2X2TS U8748 ( .A(n7440), .B(n8644), .Y(n8640) );
  NOR2XLTS U3485 ( .A(n9447), .B(n3888), .Y(n3594) );
  CLKINVX1TS U6850 ( .A(n6901), .Y(n6373) );
  AND2X2TS U2776 ( .A(n2386), .B(n9361), .Y(n2898) );
  AND2X2TS U2962 ( .A(sa10[5]), .B(n10322), .Y(n2278) );
  AND2X2TS U4846 ( .A(n4464), .B(n10084), .Y(n5006) );
  OR2X2TS U2551 ( .A(n9848), .B(n2997), .Y(n2576) );
  AND2X2TS U4449 ( .A(n10747), .B(n4282), .Y(n4734) );
  INVX1TS U4989 ( .A(n5110), .Y(n4532) );
  CLKAND2X2TS U2668 ( .A(n2940), .B(n3181), .Y(n1876) );
  NOR2XLTS U3474 ( .A(n9348), .B(n3863), .Y(n3555) );
  INVX1TS U6897 ( .A(n6640), .Y(n6914) );
  AND2X2TS U6334 ( .A(n10716), .B(n9819), .Y(n6013) );
  OR2X2TS U8763 ( .A(n8644), .B(sa20[1]), .Y(n8666) );
  AND2X2TS U4825 ( .A(n9454), .B(n3568), .Y(n4086) );
  AND2X2TS U2765 ( .A(sa21[5]), .B(n10330), .Y(n2345) );
  CLKINVX2TS U2958 ( .A(n2838), .Y(n3245) );
  NOR2XLTS U5367 ( .A(n9431), .B(n5693), .Y(n5353) );
  NAND2XLTS U1604 ( .A(n2112), .B(n2113), .Y(n1754) );
  NAND2XLTS U1592 ( .A(n2086), .B(n2087), .Y(n1716) );
  CLKINVX2TS U3125 ( .A(n2668), .Y(n3315) );
  INVX1TS U3160 ( .A(n3325), .Y(n3321) );
  CLKINVX2TS U3137 ( .A(n2167), .Y(n3026) );
  CLKAND2X2TS U2573 ( .A(n2194), .B(n2586), .Y(n2564) );
  CLKINVX2TS U8581 ( .A(n8601), .Y(n8562) );
  CLKINVX2TS U8782 ( .A(n7154), .Y(n7218) );
  CLKINVX2TS U2571 ( .A(n2586), .Y(n2036) );
  INVX1TS U2581 ( .A(n3125), .Y(n2598) );
  CLKAND2X2TS U2492 ( .A(n3130), .B(n3001), .Y(n1671) );
  CLKBUFX2TS U2545 ( .A(n2194), .Y(n2584) );
  CLKINVX2TS U4454 ( .A(n4921), .Y(n4373) );
  CLKINVX2TS U8596 ( .A(n7226), .Y(n7369) );
  CLKAND2X2TS U8524 ( .A(n8574), .B(n8579), .Y(n7358) );
  CLKINVX2TS U8766 ( .A(n8668), .Y(n8628) );
  CLKINVX2TS U6326 ( .A(n6542), .Y(n6721) );
  AND3X2TS U4459 ( .A(n9229), .B(sa33[4]), .C(n4742), .Y(n3502) );
  NAND2XLTS U8506 ( .A(n9868), .B(n9607), .Y(n8061) );
  NAND2XLTS U4124 ( .A(n4742), .B(n9229), .Y(n3844) );
  OR2X2TS U3161 ( .A(n10091), .B(n9681), .Y(n2788) );
  NOR2XLTS U7623 ( .A(sa13[3]), .B(n9570), .Y(n7753) );
  AND3X2TS U6320 ( .A(n9815), .B(n10327), .C(n6738), .Y(n6161) );
  AND2X2TS U4833 ( .A(n11190), .B(n9218), .Y(n5035) );
  OR2X2TS U2523 ( .A(n10355), .B(n9097), .Y(n2546) );
  OR2X2TS U2899 ( .A(n2848), .B(n3250), .Y(n1761) );
  OR2X2TS U6328 ( .A(n6534), .B(n9985), .Y(n6050) );
  AND2X2TS U5039 ( .A(n9193), .B(n5112), .Y(n4514) );
  NOR2XLTS U2324 ( .A(n10364), .B(n3026), .Y(n2070) );
  AND2X2TS U6928 ( .A(n6352), .B(n9452), .Y(n6316) );
  NOR3X1TS U4986 ( .A(n10313), .B(n12671), .C(n9277), .Y(n3925) );
  AND3X2TS U8354 ( .A(n10345), .B(n11181), .C(n9894), .Y(n8202) );
  OR2X2TS U8773 ( .A(n8657), .B(n9581), .Y(n7177) );
  OR2X2TS U8545 ( .A(n7369), .B(n8598), .Y(n7545) );
  NAND2XLTS U8692 ( .A(n9796), .B(n9622), .Y(n8127) );
  AND3X2TS U8136 ( .A(n8467), .B(n9585), .C(n8468), .Y(n7650) );
  OR2X2TS U2757 ( .A(n3198), .B(n9061), .Y(n1841) );
  AND2X2TS U6716 ( .A(n11202), .B(n9420), .Y(n6834) );
  OR2X2TS U2954 ( .A(n3258), .B(n9054), .Y(n1904) );
  OR2X2TS U2702 ( .A(n2924), .B(n3190), .Y(n1723) );
  NAND2XLTS U6007 ( .A(n6542), .B(n9429), .Y(n5639) );
  AND2X2TS U4423 ( .A(n9229), .B(n10367), .Y(n4280) );
  NOR2XLTS U6163 ( .A(n10710), .B(n9790), .Y(n5418) );
  NOR2XLTS U4281 ( .A(sa33[3]), .B(n9699), .Y(n3620) );
  AND2X2TS U8344 ( .A(n8414), .B(n9893), .Y(n7447) );
  AND2X2TS U3166 ( .A(n9681), .B(n10092), .Y(n3319) );
  OR2X2TS U4378 ( .A(n9698), .B(n4929), .Y(n3493) );
  NOR2XLTS U2421 ( .A(n10355), .B(n9733), .Y(n1820) );
  OR4X2TS U8322 ( .A(n9881), .B(n9593), .C(n9539), .D(sa02[2]), .Y(n7466) );
  NOR2XLTS U7707 ( .A(n10704), .B(n9580), .Y(n7784) );
  OR2X2TS U6260 ( .A(n9789), .B(n6728), .Y(n5291) );
  AND2X2TS U4638 ( .A(n11169), .B(n9211), .Y(n4977) );
  AND2X2TS U6521 ( .A(n11185), .B(n9411), .Y(n6776) );
  CLKAND2X2TS U2557 ( .A(n9062), .B(n2586), .Y(n2217) );
  AND3X2TS U8121 ( .A(n9602), .B(n9589), .C(n8463), .Y(n7691) );
  AND3X2TS U6342 ( .A(n9429), .B(sa30[4]), .C(n6542), .Y(n5300) );
  AND2X2TS U6304 ( .A(n9429), .B(n10326), .Y(n6047) );
  OR2X2TS U8588 ( .A(n8591), .B(n9570), .Y(n7249) );
  NOR2XLTS U4196 ( .A(n10309), .B(n9236), .Y(n3918) );
  OR2X2TS U3116 ( .A(n9043), .B(n9047), .Y(n2471) );
  CLKINVX1TS U4592 ( .A(n4985), .Y(n4422) );
  CLKINVX1TS U6670 ( .A(n6842), .Y(n6265) );
  CLKINVX2TS U4420 ( .A(n4938), .Y(n4783) );
  OR2X2TS U2957 ( .A(n9050), .B(n3245), .Y(n1928) );
  INVX1TS U4627 ( .A(n4980), .Y(n4982) );
  CLKINVX1TS U4787 ( .A(n5043), .Y(n4462) );
  CLKBUFX2TS U4375 ( .A(n12546), .Y(n4363) );
  OR2X2TS U2877 ( .A(n9075), .B(n3245), .Y(n1926) );
  AND2X2TS U2537 ( .A(n9062), .B(n2560), .Y(n2535) );
  INVX1TS U6705 ( .A(n6837), .Y(n6839) );
  CLKINVX2TS U8189 ( .A(n8425), .Y(n7860) );
  OR2X2TS U4447 ( .A(n9226), .B(n9925), .Y(n4283) );
  NAND2XLTS U8045 ( .A(n8425), .B(n9585), .Y(n7837) );
  CLKAND2X2TS U8157 ( .A(n8425), .B(n8477), .Y(n7847) );
  CLKAND2X2TS U8107 ( .A(n8463), .B(n8327), .Y(n7648) );
  AND3X2TS U3099 ( .A(n10091), .B(n9526), .C(n9059), .Y(n1975) );
  AND3X2TS U4438 ( .A(n9891), .B(sa33[4]), .C(n4281), .Y(n4001) );
  CLKBUFX2TS U2505 ( .A(n11452), .Y(n2042) );
  CLKINVX2TS U8195 ( .A(n8327), .Y(n7489) );
  AND3X2TS U8395 ( .A(n10730), .B(n9566), .C(n11175), .Y(n7986) );
  AND2X2TS U8367 ( .A(n9566), .B(n8539), .Y(n7455) );
  AND2X2TS U8161 ( .A(n9598), .B(n10077), .Y(n7689) );
  CLKINVX2TS U5014 ( .A(n4517), .Y(n5098) );
  OR2X2TS U2933 ( .A(n3246), .B(n9717), .Y(n2123) );
  CLKINVX2TS U6301 ( .A(n6737), .Y(n6583) );
  CLKAND2X2TS U8574 ( .A(n8590), .B(n10261), .Y(n7120) );
  CLKBUFX2TS U5023 ( .A(n12530), .Y(n4552) );
  AND3X2TS U8152 ( .A(n9854), .B(n10335), .C(n9597), .Y(n7313) );
  CLKBUFX2TS U6883 ( .A(n11723), .Y(n5983) );
  CLKBUFX2TS U3150 ( .A(n12097), .Y(n2056) );
  OR2X2TS U2901 ( .A(n9050), .B(n3237), .Y(n1947) );
  INVX1TS U2560 ( .A(n2986), .Y(n3137) );
  AND2X2TS U6842 ( .A(n9738), .B(n6674), .Y(n5575) );
  OR2X2TS U2680 ( .A(n9068), .B(n3185), .Y(n1863) );
  OR2X2TS U2704 ( .A(n9053), .B(n3177), .Y(n1884) );
  CLKBUFX2TS U6257 ( .A(n12494), .Y(n6167) );
  AND2X2TS U8727 ( .A(n9612), .B(n9560), .Y(n7418) );
  AND2X2TS U6848 ( .A(n9739), .B(n6906), .Y(n6337) );
  CLKBUFX2TS U6759 ( .A(n11759), .Y(n5744) );
  OR2X2TS U2736 ( .A(n3186), .B(n9713), .Y(n2097) );
  CLKINVX1TS U6475 ( .A(n6784), .Y(n6225) );
  INVX1TS U6510 ( .A(n6779), .Y(n6781) );
  AND2X2TS U6858 ( .A(n5753), .B(n9738), .Y(n6306) );
  AND3X2TS U8347 ( .A(n10731), .B(n11175), .C(n9535), .Y(n7969) );
  OR2X2TS U2760 ( .A(n9053), .B(n3185), .Y(n1865) );
  OR2X2TS U8364 ( .A(n9539), .B(n8491), .Y(n7465) );
  CLKINVX1TS U6900 ( .A(n6905), .Y(n6900) );
  INVX1TS U4822 ( .A(n5038), .Y(n5040) );
  CLKBUFX2TS U6932 ( .A(n10963), .Y(n5954) );
  CLKAND2X2TS U6846 ( .A(n6904), .B(n6905), .Y(n5755) );
  CLKAND2X2TS U6905 ( .A(n6904), .B(n9739), .Y(n6349) );
  OAI21X1TS U1115 ( .A0(n12667), .A1(n1258), .B0(n1259), .Y(n988) );
  NAND2XLTS U1117 ( .A(n1261), .B(n1259), .Y(n986) );
  OAI32X1TS U1120 ( .A0(n1258), .A1(n1263), .A2(n133), .B0(n1264), .B1(n1258), 
        .Y(n985) );
  OAI31X1TS U1116 ( .A0(n1260), .A1(n139), .A2(n1258), .B0(n1259), .Y(n987) );
  AND2X2TS U8590 ( .A(n9523), .B(n8590), .Y(n7253) );
  CLKBUFX2TS U6817 ( .A(n12019), .Y(n5657) );
  AND2X2TS U8714 ( .A(n9612), .B(n9505), .Y(n7438) );
  CLKBUFX2TS U4046 ( .A(n12245), .Y(n4203) );
  CLKBUFX2TS U8297 ( .A(n12635), .Y(n7992) );
  CLKBUFX2TS U2924 ( .A(n11863), .Y(n2256) );
  CLKBUFX2TS U2727 ( .A(n11887), .Y(n2323) );
  AND2X2TS U8529 ( .A(n8574), .B(n9524), .Y(n7526) );
  NAND3XLTS U7073 ( .A(n11025), .B(n10002), .C(sa20[6]), .Y(n7057) );
  CLKINVX2TS U2247 ( .A(n2612), .Y(n2012) );
  NOR2XLTS U8240 ( .A(n10732), .B(n8364), .Y(n8490) );
  AND2X2TS U8199 ( .A(n10078), .B(n9850), .Y(n7715) );
  NAND2XLTS U7960 ( .A(n11164), .B(n10749), .Y(n7582) );
  NAND2XLTS U8483 ( .A(n12076), .B(n11800), .Y(n8065) );
  CLKBUFX2TS U8486 ( .A(n11043), .Y(n7536) );
  CLKBUFX2TS U6810 ( .A(n12061), .Y(n5745) );
  NAND3XLTS U7091 ( .A(n10605), .B(n10262), .C(n11196), .Y(n7111) );
  CLKBUFX2TS U2511 ( .A(n11822), .Y(n1676) );
  CLKBUFX2TS U4403 ( .A(n11793), .Y(n4350) );
  CLKBUFX2TS U8449 ( .A(n12559), .Y(n7259) );
  CLKBUFX2TS U6418 ( .A(n12582), .Y(n5875) );
  NAND2XLTS U5660 ( .A(n11343), .B(n11695), .Y(n6009) );
  CLKBUFX2TS U8475 ( .A(n11806), .Y(n7105) );
  CLKBUFX2TS U8466 ( .A(n11082), .Y(n7550) );
  CLKBUFX2TS U6613 ( .A(n12590), .Y(n5931) );
  CLKBUFX2TS U4535 ( .A(n12586), .Y(n4075) );
  AOI22XLTS U2866 ( .A0(n12368), .A1(n11870), .B0(n11085), .B1(n11494), .Y(
        n3239) );
  NOR2XLTS U7220 ( .A(n12328), .B(n11421), .Y(n7431) );
  CLKBUFX2TS U6145 ( .A(n11752), .Y(n6287) );
  CLKBUFX2TS U2883 ( .A(n11923), .Y(n1909) );
  OR2X2TS U5876 ( .A(n11407), .B(n12505), .Y(n5700) );
  CLKBUFX2TS U8764 ( .A(n11782), .Y(n7396) );
  CLKBUFX2TS U4730 ( .A(n12579), .Y(n4131) );
  CLKBUFX2TS U2686 ( .A(n11935), .Y(n1846) );
  CLKINVX2TS U4704 ( .A(n12506), .Y(n4221) );
  OR2X2TS U5951 ( .A(n11415), .B(n12520), .Y(n5725) );
  CLKBUFX2TS U6831 ( .A(n12285), .Y(n5578) );
  OR2X2TS U6294 ( .A(n9746), .B(n6048), .Y(n6010) );
  CLKBUFX2TS U6270 ( .A(n11206), .Y(n5428) );
  OR2X2TS U6249 ( .A(n9746), .B(n6721), .Y(n6026) );
  OR2X2TS U4413 ( .A(n9656), .B(n9172), .Y(n4243) );
  NAND3XLTS U7146 ( .A(sa13[6]), .B(n10278), .C(n10261), .Y(n7248) );
  OR2X2TS U3993 ( .A(n11232), .B(n12524), .Y(n3870) );
  CLKBUFX2TS U2878 ( .A(n12603), .Y(n2247) );
  OR2X2TS U4367 ( .A(n9656), .B(n4922), .Y(n4259) );
  CLKBUFX2TS U4434 ( .A(n11785), .Y(n4351) );
  OR2X2TS U4995 ( .A(n9683), .B(n9196), .Y(n4492) );
  AND2X2TS U2501 ( .A(n9049), .B(n9051), .Y(n2559) );
  OR2X2TS U4068 ( .A(n11226), .B(n12508), .Y(n3895) );
  NAND3XLTS U7115 ( .A(n10040), .B(n10274), .C(n10001), .Y(n7176) );
  CLKBUFX2TS U6316 ( .A(n11674), .Y(n6154) );
  CLKBUFX2TS U8143 ( .A(n12369), .Y(n7682) );
  CLKBUFX2TS U2192 ( .A(n12372), .Y(n1844) );
  OAI22XLTS U5317 ( .A0(n10474), .A1(n9710), .B0(n10174), .B1(n11984), .Y(
        n5572) );
  AND2X2TS U7998 ( .A(n12162), .B(n9834), .Y(n7286) );
  NAND3BXLTS U2109 ( .AN(n9704), .B(n9725), .C(sa10[4]), .Y(n2829) );
  NOR3XLTS U5605 ( .A(n10103), .B(n11366), .C(n9755), .Y(n6102) );
  AOI31XLTS U4262 ( .A0(n11763), .A1(n12412), .A2(n10867), .B0(n11382), .Y(
        n4866) );
  NOR2XLTS U8017 ( .A(n12165), .B(n10750), .Y(n8405) );
  CLKBUFX2TS U2086 ( .A(n11566), .Y(n2252) );
  OAI22XLTS U5400 ( .A0(n12013), .A1(n10173), .B0(n10198), .B1(n11983), .Y(
        n5754) );
  NOR3XLTS U3657 ( .A(n10083), .B(n11254), .C(n9649), .Y(n4192) );
  OAI22XLTS U8469 ( .A0(n12081), .A1(n12337), .B0(n12558), .B1(n7130), .Y(
        n8575) );
  AOI22XLTS U2092 ( .A0(n10560), .A1(n10557), .B0(n11132), .B1(n9724), .Y(
        n2811) );
  OAI22XLTS U2437 ( .A0(n9931), .A1(n10016), .B0(n12555), .B1(n9928), .Y(n3104) );
  AOI22XLTS U2167 ( .A0(n10533), .A1(n10527), .B0(n11154), .B1(n9728), .Y(
        n2887) );
  NAND2XLTS U4070 ( .A(n4697), .B(n10827), .Y(n4696) );
  OAI31XLTS U5659 ( .A0(n10709), .A1(n6177), .A2(n12209), .B0(n6009), .Y(n6176) );
  NAND2XLTS U5953 ( .A(n6497), .B(n10912), .Y(n6496) );
  OAI31XLTS U3776 ( .A0(n10743), .A1(n4373), .A2(n12277), .B0(n4242), .Y(n4372) );
  AOI22XLTS U7239 ( .A0(n10305), .A1(n11505), .B0(n10311), .B1(n7467), .Y(
        n7464) );
  AOI31XLTS U7364 ( .A0(n11528), .A1(n11921), .A2(n10338), .B0(n10706), .Y(
        n7718) );
  OAI21XLTS U2142 ( .A0(n10560), .A1(n12301), .B0(n11869), .Y(n2862) );
  NOR3XLTS U5577 ( .A(n10075), .B(n11360), .C(n9751), .Y(n6058) );
  NAND2XLTS U6113 ( .A(n6639), .B(n10550), .Y(n6638) );
  NAND3XLTS U8002 ( .A(n11890), .B(n11645), .C(n9527), .Y(n7300) );
  OAI22XLTS U8234 ( .A0(n10093), .A1(n9528), .B0(n10744), .B1(n9833), .Y(n8486) );
  CLKBUFX2TS U8348 ( .A(n11890), .Y(n7458) );
  NAND3BXLTS U2184 ( .AN(n9708), .B(n9729), .C(n10727), .Y(n2905) );
  NOR3XLTS U3629 ( .A(n10055), .B(n11261), .C(n9645), .Y(n4148) );
  NAND2XLTS U3995 ( .A(n4625), .B(n10854), .Y(n4624) );
  CLKBUFX2TS U2161 ( .A(n11577), .Y(n2319) );
  OAI22XLTS U7447 ( .A0(n11103), .A1(n9845), .B0(n10061), .B1(n10717), .Y(
        n7839) );
  NAND2XLTS U5878 ( .A(n6425), .B(n10884), .Y(n6424) );
  OR2X2TS U6458 ( .A(n12220), .B(n10908), .Y(n5450) );
  CLKBUFX2TS U4844 ( .A(n10804), .Y(n4130) );
  NAND2XLTS U2272 ( .A(n12555), .B(n10685), .Y(n2984) );
  CLKBUFX2TS U4368 ( .A(n12275), .Y(n3841) );
  CLKBUFX2TS U2936 ( .A(n11875), .Y(n2457) );
  CLKBUFX2TS U6532 ( .A(n10908), .Y(n5874) );
  CLKBUFX2TS U6343 ( .A(n11671), .Y(n6025) );
  AOI22XLTS U2859 ( .A0(n11115), .A1(n1758), .B0(n12132), .B1(n9975), .Y(n3233) );
  NAND2XLTS U6000 ( .A(n12211), .B(n9766), .Y(n6046) );
  OR2X2TS U6653 ( .A(n12243), .B(n10937), .Y(n5516) );
  CLKBUFX2TS U8495 ( .A(n11849), .Y(n8093) );
  NAND2XLTS U8628 ( .A(n11837), .B(n12068), .Y(n7394) );
  NOR2XLTS U2826 ( .A(n10556), .B(n10578), .Y(n3225) );
  OAI21XLTS U4791 ( .A0(n11285), .A1(n12051), .B0(n11280), .Y(n5050) );
  OR2X2TS U2690 ( .A(n10532), .B(n11577), .Y(n1886) );
  OAI21XLTS U4596 ( .A0(n11334), .A1(n12060), .B0(n11326), .Y(n4992) );
  CLKBUFX2TS U2739 ( .A(n11899), .Y(n2413) );
  OAI22XLTS U7451 ( .A0(n10286), .A1(n11610), .B0(n10712), .B1(n10718), .Y(
        n7858) );
  NAND2XLTS U8110 ( .A(n10337), .B(n10657), .Y(n7663) );
  CLKBUFX2TS U4408 ( .A(n10129), .Y(n3486) );
  NAND2XLTS U4117 ( .A(n12275), .B(n9929), .Y(n4279) );
  CLKBUFX2TS U4389 ( .A(n11416), .Y(n3630) );
  OAI21XLTS U6674 ( .A0(n11319), .A1(n11972), .B0(n11323), .Y(n6849) );
  OR2X2TS U4575 ( .A(n12270), .B(n10831), .Y(n3695) );
  CLKBUFX2TS U8686 ( .A(n11831), .Y(n8159) );
  CLKBUFX2TS U4732 ( .A(n10827), .Y(n4119) );
  OAI21XLTS U6479 ( .A0(n11271), .A1(n11975), .B0(n11277), .Y(n6791) );
  OR2X2TS U4770 ( .A(n12246), .B(n4130), .Y(n3761) );
  CLKBUFX2TS U8089 ( .A(n11903), .Y(n7724) );
  CLKBUFX2TS U2453 ( .A(n12554), .Y(n2562) );
  CLKBUFX2TS U8759 ( .A(n12107), .Y(n7066) );
  OR2X2TS U2887 ( .A(n10561), .B(n2252), .Y(n1949) );
  AND2X2TS U8092 ( .A(n11522), .B(n10285), .Y(n7692) );
  OAI31XLTS U1721 ( .A0(n2341), .A1(n9069), .A2(n10543), .B0(n2343), .Y(n2331)
         );
  CLKBUFX2TS U4987 ( .A(n11713), .Y(n4482) );
  AOI31XLTS U7491 ( .A0(n12101), .A1(n12119), .A2(n12334), .B0(n10627), .Y(
        n7899) );
  OAI22XLTS U5597 ( .A0(n10568), .A1(n10462), .B0(n10525), .B1(n12026), .Y(
        n6093) );
  AOI32XLTS U2174 ( .A0(n10727), .A1(n2898), .A2(n11490), .B0(n9944), .B1(
        n9988), .Y(n2896) );
  INVX1TS U1978 ( .A(n2306), .Y(n2093) );
  CLKBUFX2TS U8659 ( .A(n11776), .Y(n7157) );
  OAI31XLTS U6357 ( .A0(sa12[2]), .A1(n9436), .A2(n12415), .B0(n6431), .Y(
        n6745) );
  CLKBUFX2TS U4896 ( .A(n12493), .Y(n4575) );
  INVXLTS U2631 ( .A(n2346), .Y(n3163) );
  NAND2XLTS U4326 ( .A(n4903), .B(n10159), .Y(n4902) );
  CLKBUFX2TS U8108 ( .A(n12355), .Y(n7733) );
  NOR2XLTS U7413 ( .A(n11796), .B(n11425), .Y(n7796) );
  NOR3XLTS U8648 ( .A(n10705), .B(n11776), .C(n8628), .Y(n8635) );
  AOI31XLTS U7534 ( .A0(n11795), .A1(n11836), .A2(n12148), .B0(n10617), .Y(
        n7946) );
  OAI22XLTS U8699 ( .A0(n11603), .A1(n11830), .B0(n11776), .B1(n11419), .Y(
        n8654) );
  AOI22XLTS U5288 ( .A0(n10909), .A1(n12510), .B0(n9635), .B1(n11276), .Y(
        n5488) );
  CLKINVX2TS U6798 ( .A(n5955), .Y(n6298) );
  CLKBUFX2TS U8098 ( .A(n12633), .Y(n7325) );
  CLKBUFX2TS U6494 ( .A(n12513), .Y(n5866) );
  NOR2XLTS U8127 ( .A(n9861), .B(n11611), .Y(n8316) );
  OAI211XLTS U2652 ( .A0(n2692), .A1(n10672), .B0(n2879), .C0(n2902), .Y(n3176) );
  AOI22XLTS U3417 ( .A0(n10832), .A1(n12514), .B0(n9636), .B1(n11327), .Y(
        n3733) );
  INVX1TS U6794 ( .A(n6630), .Y(n6890) );
  CLKBUFX2TS U4939 ( .A(n12541), .Y(n4506) );
  NAND2XLTS U6208 ( .A(n6702), .B(n10141), .Y(n6701) );
  OAI32X1TS U5952 ( .A0(sa23[6]), .A1(n9754), .A2(n11311), .B0(n6496), .B1(
        n10104), .Y(n5385) );
  AOI31XLTS U5399 ( .A0(n9345), .A1(n5753), .A2(n5954), .B0(n5754), .Y(n5752)
         );
  AOI22XLTS U1992 ( .A0(n10564), .A1(n12603), .B0(n9971), .B1(n11130), .Y(
        n2712) );
  AOI22XLTS U1993 ( .A0(n9972), .A1(n11923), .B0(n10248), .B1(n11496), .Y(
        n2711) );
  INVXLTS U2828 ( .A(n2279), .Y(n3223) );
  OAI31XLTS U4474 ( .A0(n11168), .A1(n9240), .A2(n12403), .B0(n4631), .Y(n4946) );
  CLKBUFX2TS U8473 ( .A(n12094), .Y(n7229) );
  CLKBUFX2TS U2455 ( .A(n11911), .Y(n2040) );
  INVX1TS U2020 ( .A(n2239), .Y(n2119) );
  NOR2XLTS U7390 ( .A(n12102), .B(n12081), .Y(n7764) );
  OAI22XLTS U3677 ( .A0(n10372), .A1(n10438), .B0(n10387), .B1(n11994), .Y(
        n4227) );
  OAI31XLTS U1686 ( .A0(n2274), .A1(n9075), .A2(n10569), .B0(n2276), .Y(n2264)
         );
  CLKBUFX2TS U4611 ( .A(n12517), .Y(n4066) );
  AND2X2TS U7549 ( .A(n9878), .B(n11119), .Y(n7293) );
  OAI32X1TS U5877 ( .A0(sa12[6]), .A1(n9750), .A2(n11263), .B0(n6424), .B1(
        n10076), .Y(n5346) );
  NOR3XLTS U8462 ( .A(n10738), .B(n12096), .C(n8562), .Y(n8569) );
  AOI31XLTS U7311 ( .A0(n9535), .A1(n10643), .A2(n9539), .B0(n7621), .Y(n7618)
         );
  OAI22XLTS U5625 ( .A0(n10573), .A1(n10469), .B0(n10535), .B1(n12041), .Y(
        n6137) );
  OAI22XLTS U3649 ( .A0(n10378), .A1(n10446), .B0(n10399), .B1(n12009), .Y(
        n4183) );
  AOI31XLTS U7667 ( .A0(n12094), .A1(n11849), .A2(n12560), .B0(n11874), .Y(
        n8082) );
  CLKBUFX2TS U8334 ( .A(n11118), .Y(n8209) );
  OAI21XLTS U7665 ( .A0(n11563), .A1(n10733), .B0(n11457), .Y(n8085) );
  AOI31XLTS U8030 ( .A0(sa02[7]), .A1(n8414), .A2(n10305), .B0(n8415), .Y(
        n8409) );
  AOI21XLTS U8025 ( .A0(n12156), .A1(n10097), .B0(n7629), .Y(n8412) );
  OAI32X1TS U4069 ( .A0(sa22[6]), .A1(n9648), .A2(n11292), .B0(n4696), .B1(
        n10084), .Y(n3587) );
  CLKINVX2TS U8325 ( .A(n8385), .Y(n8408) );
  OAI211XLTS U2849 ( .A0(n2725), .A1(n10659), .B0(n2803), .C0(n2826), .Y(n3236) );
  AOI22XLTS U1869 ( .A0(n9048), .A1(n10583), .B0(n11454), .B1(n11005), .Y(
        n2574) );
  AOI22XLTS U5313 ( .A0(n10936), .A1(n12526), .B0(n9633), .B1(n11324), .Y(
        n5554) );
  AOI31XLTS U7752 ( .A0(n11777), .A1(n11831), .A2(n12329), .B0(n11541), .Y(
        n8148) );
  AOI22XLTS U3442 ( .A0(n10805), .A1(n12498), .B0(n9638), .B1(n11279), .Y(
        n3799) );
  NAND3XLTS U8654 ( .A(n9506), .B(n11059), .C(n8644), .Y(n7428) );
  INVX1TS U7733 ( .A(n7798), .Y(n7429) );
  AOI211XLTS U1610 ( .A0(n10700), .A1(n2822), .B0(n12125), .C0(n2126), .Y(
        n2116) );
  AOI32XLTS U2099 ( .A0(n10699), .A1(n2822), .A2(n11496), .B0(n9947), .B1(
        n9976), .Y(n2820) );
  CLKBUFX2TS U6689 ( .A(n12529), .Y(n5922) );
  CLKBUFX2TS U4806 ( .A(n12500), .Y(n4122) );
  CLKINVX2TS U6856 ( .A(n5586), .Y(n6297) );
  NOR2X1TS U5382 ( .A(n11972), .B(n12272), .Y(n5722) );
  NAND2XLTS U2424 ( .A(n9062), .B(n10610), .Y(n3099) );
  NOR2X1TS U3488 ( .A(n12051), .B(n12214), .Y(n3892) );
  OAI22XLTS U2309 ( .A0(n12555), .A1(n10304), .B0(n9720), .B1(n10603), .Y(
        n3013) );
  AND2X2TS U4729 ( .A(n9150), .B(n10895), .Y(n3793) );
  OAI22XLTS U2307 ( .A0(n1807), .A1(n12161), .B0(n2607), .B1(n10603), .Y(n3014) );
  OAI32X1TS U8480 ( .A0(n11196), .A1(n7547), .A2(n11044), .B0(n8582), .B1(
        n11197), .Y(n7743) );
  OAI21XLTS U3694 ( .A0(n10742), .A1(n9652), .B0(n12283), .Y(n4017) );
  OAI22XLTS U2305 ( .A0(n2014), .A1(n11588), .B0(n9721), .B1(n11045), .Y(n3015) );
  AOI22XLTS U2986 ( .A0(n10966), .A1(n11538), .B0(n12110), .B1(n11067), .Y(
        n3268) );
  NOR3XLTS U2790 ( .A(sa10[2]), .B(n9076), .C(n11881), .Y(n3206) );
  NAND2XLTS U8042 ( .A(n9897), .B(n12142), .Y(n8424) );
  OAI22XLTS U4032 ( .A0(n4121), .A1(n11290), .B0(n4660), .B1(n9161), .Y(n4658)
         );
  CLKINVX2TS U2294 ( .A(n2518), .Y(n1662) );
  OAI31XLTS U3925 ( .A0(n9200), .A1(n4515), .A2(n4807), .B0(n4547), .Y(n4538)
         );
  OAI22XLTS U7918 ( .A0(n10065), .A1(n9862), .B0(n10074), .B1(n11557), .Y(
        n8318) );
  CLKBUFX2TS U4579 ( .A(n12222), .Y(n3701) );
  OAI22XLTS U2230 ( .A0(n9999), .A1(n9931), .B0(n10695), .B1(n10684), .Y(n2948) );
  NOR2XLTS U3922 ( .A(n10407), .B(n11713), .Y(n4543) );
  AOI22XLTS U5543 ( .A0(n11395), .A1(n10496), .B0(n9990), .B1(n11668), .Y(
        n6008) );
  OAI21XLTS U7189 ( .A0(n12307), .A1(n7369), .B0(n7370), .Y(n7361) );
  OAI22XLTS U7629 ( .A0(n12103), .A1(n10627), .B0(n10328), .B1(n11849), .Y(
        n8051) );
  OAI22XLTS U7148 ( .A0(n7252), .A1(n11808), .B0(n10021), .B1(n11802), .Y(
        n7251) );
  OAI21XLTS U5546 ( .A0(sa30[3]), .A1(n9742), .B0(n12204), .Y(n5803) );
  OAI22XLTS U3957 ( .A0(n4065), .A1(n11338), .B0(n4588), .B1(n9153), .Y(n4586)
         );
  OAI22XLTS U7507 ( .A0(n9809), .A1(n10600), .B0(n11843), .B1(n12150), .Y(
        n7912) );
  OAI22XLTS U2813 ( .A0(n2244), .A1(n11883), .B0(n11876), .B1(n11864), .Y(
        n3214) );
  OAI22XLTS U5840 ( .A0(n5865), .A1(n11263), .B0(n6388), .B1(n9359), .Y(n6386)
         );
  AOI21XLTS U1999 ( .A0(n10654), .A1(n10243), .B0(n11430), .Y(n2715) );
  NOR2X1TS U5370 ( .A(n11975), .B(n12264), .Y(n5697) );
  AND2X2TS U4534 ( .A(n9138), .B(n10911), .Y(n3727) );
  OAI22XLTS U5559 ( .A0(n5410), .A1(n10416), .B0(n12203), .B1(n11671), .Y(
        n6032) );
  NAND2XLTS U5804 ( .A(n12293), .B(n10249), .Y(n6348) );
  NAND3XLTS U1938 ( .A(n2668), .B(n9955), .C(n10096), .Y(n2667) );
  OAI22XLTS U1773 ( .A0(n2423), .A1(n11470), .B0(n2239), .B1(n11864), .Y(n2421) );
  OAI22XLTS U1518 ( .A0(n9979), .A1(n11882), .B0(n10640), .B1(n10256), .Y(
        n1906) );
  OAI22XLTS U2035 ( .A0(n11063), .A1(n11458), .B0(n9046), .B1(n9924), .Y(n2746) );
  OAI22XLTS U1776 ( .A0(n2431), .A1(n11120), .B0(n10570), .B1(n10256), .Y(
        n2426) );
  NOR2XLTS U1778 ( .A(n10243), .B(n11472), .Y(n2425) );
  OAI22XLTS U5915 ( .A0(n5921), .A1(n11311), .B0(n6460), .B1(n9367), .Y(n6458)
         );
  AOI22XLTS U7666 ( .A0(n11570), .A1(n11445), .B0(n11627), .B1(n10687), .Y(
        n8084) );
  OAI22XLTS U7325 ( .A0(n10285), .A1(n11557), .B0(n11528), .B1(n10707), .Y(
        n7657) );
  OAI32X1TS U6207 ( .A0(n10044), .A1(n11401), .A2(n9985), .B0(n6701), .B1(
        sa30[6]), .Y(n6175) );
  OAI22XLTS U1749 ( .A0(n2387), .A1(n11141), .B0(n10543), .B1(n10280), .Y(
        n2382) );
  NOR2XLTS U1751 ( .A(n10267), .B(n11484), .Y(n2381) );
  INVX1TS U8684 ( .A(n7426), .Y(n7920) );
  OAI32X1TS U8665 ( .A0(sa20[6]), .A1(n7404), .A2(n10600), .B0(n8646), .B1(
        n10040), .Y(n7774) );
  AND2X2TS U6612 ( .A(n9349), .B(n10874), .Y(n5548) );
  OAI22XLTS U7620 ( .A0(n12114), .A1(n12336), .B0(n11933), .B1(n11113), .Y(
        n8049) );
  OAI21XLTS U8246 ( .A0(n10085), .A1(n11645), .B0(n8358), .Y(n8495) );
  AOI31XLTS U8646 ( .A0(sa20[4]), .A1(n9612), .A2(n11784), .B0(n7430), .Y(
        n8636) );
  OAI22XLTS U5639 ( .A0(n5315), .A1(n9356), .B0(n5639), .B1(n11401), .Y(n6148)
         );
  OAI22XLTS U8643 ( .A0(n11468), .A1(n12329), .B0(n11838), .B1(n11420), .Y(
        n8639) );
  AND2X2TS U6021 ( .A(n9356), .B(n10412), .Y(n5302) );
  CLKBUFX2TS U4900 ( .A(n10802), .Y(n3668) );
  AOI22XLTS U6019 ( .A0(n12449), .A1(n9989), .B0(n11379), .B1(n10563), .Y(
        n6555) );
  INVX1TS U6034 ( .A(n5809), .Y(n6011) );
  CLKBUFX2TS U6066 ( .A(n10241), .Y(n5797) );
  AOI21XLTS U7912 ( .A0(n10065), .A1(n9551), .B0(n11509), .Y(n8310) );
  AND2X2TS U6417 ( .A(n9334), .B(n10858), .Y(n5482) );
  NAND2XLTS U4233 ( .A(n4840), .B(n10148), .Y(n4839) );
  OAI22XLTS U7533 ( .A0(n11842), .A1(n12327), .B0(n10293), .B1(n12067), .Y(
        n7947) );
  OAI22XLTS U1746 ( .A0(n2379), .A1(n11482), .B0(n2306), .B1(n11887), .Y(n2377) );
  OAI32X1TS U4325 ( .A0(n10748), .A1(n11707), .A2(n9925), .B0(n4902), .B1(
        sa33[6]), .Y(n4371) );
  AOI22XLTS U4136 ( .A0(n12377), .A1(n9933), .B0(n10784), .B1(n10380), .Y(
        n4755) );
  AOI32XLTS U7517 ( .A0(n7180), .A1(n7421), .A2(n11765), .B0(n11795), .B1(
        n7421), .Y(n7926) );
  OAI22XLTS U7766 ( .A0(n7802), .A1(n12069), .B0(n7071), .B1(n9802), .Y(n8160)
         );
  CLKBUFX2TS U4183 ( .A(n10125), .Y(n3984) );
  OAI22XLTS U5257 ( .A0(n5410), .A1(n12196), .B0(n5411), .B1(n11672), .Y(n5409) );
  NAND2XLTS U2488 ( .A(n12554), .B(n11638), .Y(n3127) );
  OAI22XLTS U7415 ( .A0(n11820), .A1(n12330), .B0(n11539), .B1(n12150), .Y(
        n7792) );
  OAI22XLTS U3375 ( .A0(n3612), .A1(n12066), .B0(n3613), .B1(n11386), .Y(n3611) );
  AOI31XLTS U8460 ( .A0(sa13[4]), .A1(n8574), .A2(n11451), .B0(n7514), .Y(
        n8570) );
  OAI22XLTS U7489 ( .A0(n11485), .A1(n10682), .B0(n11872), .B1(n11848), .Y(
        n7901) );
  OAI22XLTS U7490 ( .A0(n12319), .A1(n12558), .B0(n10677), .B1(n12304), .Y(
        n7900) );
  OAI22XLTS U1494 ( .A0(n9991), .A1(n11905), .B0(n10649), .B1(n10280), .Y(
        n1843) );
  NOR2X1TS U5247 ( .A(n12241), .B(n12410), .Y(n5380) );
  OAI31XLTS U2145 ( .A0(n9936), .A1(n9281), .A2(n11466), .B0(n2867), .Y(n2865)
         );
  CLKBUFX2TS U3051 ( .A(n12110), .Y(n2628) );
  OAI31XLTS U2220 ( .A0(n9940), .A1(n9361), .A2(n11478), .B0(n2943), .Y(n2941)
         );
  OAI22XLTS U2157 ( .A0(n2881), .A1(n11631), .B0(n11434), .B1(n10279), .Y(
        n2876) );
  NOR2X1TS U3365 ( .A(n12244), .B(n12422), .Y(n3582) );
  OAI22XLTS U2158 ( .A0(n11583), .A1(n10268), .B0(n9991), .B1(n11630), .Y(
        n2875) );
  INVX1TS U3138 ( .A(n2777), .Y(n2514) );
  AOI32XLTS U5647 ( .A0(n5625), .A1(n11670), .A2(sa30[4]), .B0(n10241), .B1(
        n11668), .Y(n6160) );
  OAI22XLTS U2246 ( .A0(n2617), .A1(n12565), .B0(n2012), .B1(n10684), .Y(n2958) );
  AND2X2TS U8300 ( .A(n10356), .B(n9833), .Y(n7608) );
  NAND2XLTS U8292 ( .A(sa02[4]), .B(n12177), .Y(n8522) );
  NOR2X1TS U5236 ( .A(n12218), .B(n12394), .Y(n5341) );
  NOR2XLTS U7452 ( .A(n12488), .B(n12142), .Y(n7854) );
  AOI21XLTS U1957 ( .A0(n10667), .A1(n10267), .B0(n11436), .Y(n2682) );
  NOR2X1TS U3354 ( .A(n12268), .B(n12438), .Y(n3543) );
  OAI22XLTS U2083 ( .A0(n11572), .A1(n10244), .B0(n9979), .B1(n11612), .Y(
        n2799) );
  OAI22XLTS U3756 ( .A0(n3517), .A1(n9169), .B0(n3844), .B1(n11707), .Y(n4345)
         );
  OAI22XLTS U2082 ( .A0(n2805), .A1(n11613), .B0(n11428), .B1(n10255), .Y(
        n2800) );
  AOI22XLTS U6775 ( .A0(n9973), .A1(n5955), .B0(n12300), .B1(n5586), .Y(n6881)
         );
  AND2X2TS U4982 ( .A(n9678), .B(n9901), .Y(n3636) );
  NAND2XLTS U6789 ( .A(n12293), .B(n10177), .Y(n6888) );
  OAI22XLTS U8457 ( .A0(n11486), .A1(n12560), .B0(n12121), .B1(n11801), .Y(
        n8573) );
  OAI22XLTS U8709 ( .A0(n7191), .A1(n9809), .B0(n11776), .B1(n11467), .Y(n8662) );
  AOI32XLTS U7474 ( .A0(n7252), .A1(n7531), .A2(n12077), .B0(n12100), .B1(
        n7531), .Y(n7879) );
  AOI32XLTS U4022 ( .A0(sa11[4]), .A1(n10907), .A2(n4061), .B0(n10405), .B1(
        n10905), .Y(n4649) );
  OAI22XLTS U3574 ( .A0(n10425), .A1(n10844), .B0(n11412), .B1(n12403), .Y(
        n4062) );
  OAI31XLTS U4110 ( .A0(n9892), .A1(n9225), .A2(n12064), .B0(n4369), .Y(n4729)
         );
  OAI22XLTS U5457 ( .A0(n10506), .A1(n10896), .B0(n11204), .B1(n12418), .Y(
        n5862) );
  AOI21XLTS U4154 ( .A0(n10759), .A1(n12276), .B0(n11709), .Y(n4773) );
  OAI211XLTS U4788 ( .A0(n10815), .A1(n9912), .B0(n5050), .C0(n4675), .Y(n5048) );
  NOR2XLTS U4156 ( .A(n12389), .B(n11707), .Y(n4774) );
  AOI31XLTS U5902 ( .A0(n6063), .A1(n10072), .A2(n10162), .B0(n6215), .Y(n6447) );
  AOI32XLTS U5905 ( .A0(n9435), .A1(n10862), .A2(n5861), .B0(n10581), .B1(
        n10862), .Y(n6449) );
  OAI22XLTS U6369 ( .A0(n5865), .A1(n10209), .B0(n5831), .B1(n12025), .Y(n6755) );
  AOI21XLTS U6037 ( .A0(n10985), .A1(n12210), .B0(n11403), .Y(n6573) );
  OR2X2TS U6041 ( .A(n11677), .B(n9993), .Y(n5806) );
  NOR2XLTS U6039 ( .A(n12441), .B(n11401), .Y(n6574) );
  OAI22XLTS U5281 ( .A0(n5477), .A1(n11265), .B0(n5348), .B1(n10461), .Y(n5476) );
  AOI22XLTS U5287 ( .A0(n11693), .A1(n11973), .B0(n12224), .B1(n12263), .Y(
        n5489) );
  NAND2XLTS U4776 ( .A(n10381), .B(n10471), .Y(n4223) );
  OR2X2TS U4158 ( .A(n11791), .B(n10121), .Y(n4020) );
  AND2X2TS U6769 ( .A(n11019), .B(n11991), .Y(n6341) );
  AND2X2TS U4138 ( .A(n9169), .B(n10163), .Y(n3504) );
  OR2X2TS U8673 ( .A(n11065), .B(n10673), .Y(n7209) );
  AOI22XLTS U3416 ( .A0(n11738), .A1(n12057), .B0(n12259), .B1(n12221), .Y(
        n3734) );
  OAI22XLTS U3544 ( .A0(n10759), .A1(n9919), .B0(n10152), .B1(n12066), .Y(
        n4011) );
  OAI22XLTS U3410 ( .A0(n3722), .A1(n11340), .B0(n3550), .B1(n10447), .Y(n3721) );
  AOI22XLTS U4920 ( .A0(n10137), .A1(n12619), .B0(n10812), .B1(n11701), .Y(
        n5099) );
  OAI22XLTS U5420 ( .A0(n10985), .A1(n9941), .B0(n10150), .B1(n12197), .Y(
        n5795) );
  AOI31XLTS U4019 ( .A0(n4153), .A1(n10052), .A2(n10136), .B0(n4412), .Y(n4647) );
  AOI31XLTS U3938 ( .A0(n9204), .A1(n10410), .A2(n10307), .B0(n4572), .Y(n4557) );
  OAI211XLTS U5802 ( .A0(n11991), .A1(n5578), .B0(n6348), .C0(n5966), .Y(n6347) );
  AOI31XLTS U5805 ( .A0(n9782), .A1(n11748), .A2(n10197), .B0(n11736), .Y(
        n6346) );
  AOI22XLTS U5819 ( .A0(n11355), .A1(n11759), .B0(n10947), .B1(n10201), .Y(
        n6366) );
  OAI22XLTS U5816 ( .A0(n5662), .A1(n10225), .B0(n11020), .B1(n12286), .Y(
        n6371) );
  AOI31XLTS U3926 ( .A0(n9921), .A1(n12568), .A2(n10111), .B0(n12530), .Y(
        n4537) );
  OAI31XLTS U2121 ( .A0(n10028), .A1(n9716), .A2(n12347), .B0(n2843), .Y(n2842) );
  OAI32XLTS U3924 ( .A0(n12380), .A1(n9193), .A2(n9197), .B0(n10791), .B1(
        n12379), .Y(n4539) );
  OAI31XLTS U2289 ( .A0(n2998), .A1(n12679), .A2(n10291), .B0(n1665), .Y(n2969) );
  OAI21XLTS U3936 ( .A0(n10796), .A1(n9190), .B0(n9175), .Y(n4563) );
  OAI22XLTS U3934 ( .A0(n10791), .A1(n12540), .B0(n12413), .B1(n12531), .Y(
        n4567) );
  NAND3XLTS U4274 ( .A(n4876), .B(n4841), .C(sa00[4]), .Y(n4869) );
  OAI31XLTS U2196 ( .A0(n10060), .A1(n9712), .A2(n1884), .B0(n2919), .Y(n2918)
         );
  NAND4XLTS U7662 ( .A(n8084), .B(n8085), .C(n7768), .D(n7754), .Y(n8083) );
  AOI211XLTS U1517 ( .A0(n11930), .A1(n10259), .B0(n1905), .C0(n1906), .Y(
        n1902) );
  OAI211XLTS U3690 ( .A0(n12276), .A1(n3493), .B0(n4241), .C0(n4242), .Y(n4240) );
  AOI31XLTS U7269 ( .A0(n9523), .A1(n10278), .A2(n7528), .B0(n7529), .Y(n7521)
         );
  OAI22XLTS U2080 ( .A0(n11571), .A1(n12466), .B0(n10574), .B1(n9079), .Y(
        n2804) );
  OAI22XLTS U4486 ( .A0(n4065), .A1(n10105), .B0(n4031), .B1(n12008), .Y(n4956) );
  NOR2XLTS U1685 ( .A(n12461), .B(n12347), .Y(n2269) );
  OAI22XLTS U1683 ( .A0(n12167), .A1(n10993), .B0(n9980), .B1(n10659), .Y(
        n2271) );
  OAI22XLTS U3705 ( .A0(n10757), .A1(n9913), .B0(n10503), .B1(n10765), .Y(
        n4269) );
  OAI22XLTS U2051 ( .A0(n2769), .A1(n11015), .B0(n10524), .B1(n10629), .Y(
        n2768) );
  NAND4XLTS U7436 ( .A(n7828), .B(n7829), .C(n11597), .D(n11509), .Y(n7810) );
  INVXLTS U3042 ( .A(n3071), .Y(n3293) );
  NOR2XLTS U7830 ( .A(n12172), .B(n11587), .Y(n8238) );
  OAI31XLTS U7853 ( .A0(sa02[3]), .A1(n11952), .A2(n8237), .B0(n8261), .Y(
        n8242) );
  OAI22XLTS U5642 ( .A0(n9743), .A1(n9759), .B0(n9763), .B1(n9941), .Y(n6152)
         );
  OAI22XLTS U3911 ( .A0(n10790), .A1(n11380), .B0(n9901), .B1(n11714), .Y(
        n4531) );
  OAI22XLTS U7801 ( .A0(n10347), .A1(n10098), .B0(n11188), .B1(n11646), .Y(
        n8198) );
  OAI22XLTS U5793 ( .A0(n11020), .A1(n9982), .B0(n6320), .B1(n11752), .Y(n6333) );
  OAI22XLTS U3759 ( .A0(n9653), .A1(n9661), .B0(n9665), .B1(n9919), .Y(n4349)
         );
  OAI211XLTS U6102 ( .A0(n12286), .A1(n11371), .B0(n6630), .C0(n6278), .Y(
        n6629) );
  AOI22XLTS U7844 ( .A0(n8180), .A1(n10642), .B0(n10089), .B1(n11503), .Y(
        n8255) );
  AOI33X1TS U7864 ( .A0(n8271), .A1(n10090), .A2(n10345), .B0(n8272), .B1(
        n10642), .B2(sa02[2]), .Y(n8266) );
  AOI31XLTS U7560 ( .A0(n10093), .A1(n10347), .A2(n12162), .B0(n11575), .Y(
        n7985) );
  OAI31XLTS U3105 ( .A0(n9522), .A1(n9070), .A2(n11531), .B0(n1967), .Y(n3320)
         );
  AOI22XLTS U7307 ( .A0(n10333), .A1(n7610), .B0(n12179), .B1(n7296), .Y(n7602) );
  AOI22XLTS U7305 ( .A0(n11910), .A1(n9481), .B0(n12479), .B1(n7467), .Y(n7604) );
  AOI22XLTS U7304 ( .A0(n11134), .A1(n7593), .B0(n10310), .B1(n11498), .Y(
        n7605) );
  OAI21XLTS U1927 ( .A0(n9042), .A1(n2652), .B0(n12118), .Y(n2493) );
  OAI22XLTS U1669 ( .A0(n2239), .A1(n12461), .B0(n10574), .B1(n10999), .Y(
        n2238) );
  OAI32XLTS U5807 ( .A0(n12012), .A1(n6351), .A2(n6352), .B0(n11019), .B1(
        n12011), .Y(n6350) );
  OAI22XLTS U3000 ( .A0(n2761), .A1(n11858), .B0(n2153), .B1(n10624), .Y(n3274) );
  OAI22XLTS U7633 ( .A0(n7123), .A1(n11128), .B0(n12114), .B1(n10021), .Y(
        n8059) );
  AOI22XLTS U1904 ( .A0(n11823), .A1(n11513), .B0(n12091), .B1(n2619), .Y(
        n2618) );
  OAI22XLTS U7704 ( .A0(n11818), .A1(n12149), .B0(n11605), .B1(n11070), .Y(
        n8115) );
  OAI31XLTS U2990 ( .A0(sa03[2]), .A1(n11853), .A2(n9952), .B0(n2143), .Y(
        n3269) );
  OAI32X1TS U8041 ( .A0(n10341), .A1(n7727), .A2(n11559), .B0(n8424), .B1(
        n10340), .Y(n8031) );
  OR2X2TS U8698 ( .A(n11939), .B(n9576), .Y(n7067) );
  AOI31XLTS U8572 ( .A0(n8603), .A1(n9864), .A2(n10277), .B0(n8048), .Y(n8612)
         );
  OAI21XLTS U1461 ( .A0(sa10[7]), .A1(n9119), .B0(n12459), .Y(n1768) );
  OAI22XLTS U1500 ( .A0(n11619), .A1(n11626), .B0(n11142), .B1(n11630), .Y(
        n1856) );
  OAI22XLTS U2155 ( .A0(n11582), .A1(n12482), .B0(n10547), .B1(n9072), .Y(
        n2880) );
  AOI22XLTS U7198 ( .A0(n11059), .A1(n10670), .B0(n10289), .B1(n7215), .Y(
        n7388) );
  NOR2XLTS U1720 ( .A(n12475), .B(n12354), .Y(n2336) );
  OAI22XLTS U1718 ( .A0(n12173), .A1(n10977), .B0(n9992), .B1(n10672), .Y(
        n2338) );
  AOI32XLTS U8238 ( .A0(n10744), .A1(n8261), .A2(n11639), .B0(n11187), .B1(
        n8261), .Y(n8489) );
  OAI31XLTS U7196 ( .A0(n10036), .A1(n9496), .A2(n11766), .B0(n7385), .Y(n7383) );
  AOI22XLTS U7402 ( .A0(n11783), .A1(n10613), .B0(n11053), .B1(n7784), .Y(
        n7783) );
  OAI21XLTS U1448 ( .A0(sa21[7]), .A1(n9123), .B0(n12476), .Y(n1730) );
  AOI31XLTS U8458 ( .A0(n10262), .A1(n11197), .A2(n11629), .B0(n7142), .Y(
        n8571) );
  OAI31XLTS U7478 ( .A0(n11934), .A1(n9867), .A2(n9841), .B0(n7563), .Y(n7881)
         );
  AND2X2TS U2266 ( .A(n10689), .B(n9963), .Y(n2202) );
  AOI221XLTS U5835 ( .A0(n5333), .A1(n9380), .B0(n11682), .B1(n11973), .C0(
        n6383), .Y(n6382) );
  OAI22XLTS U7506 ( .A0(n11764), .A1(n11071), .B0(n7080), .B1(n10665), .Y(
        n7913) );
  INVX1TS U7695 ( .A(n8057), .Y(n8096) );
  OAI32XLTS U2234 ( .A0(n12159), .A1(n10350), .A2(n2036), .B0(n10012), .B1(
        n11948), .Y(n2953) );
  CLKINVX2TS U2465 ( .A(n2201), .Y(n2587) );
  OAI22XLTS U7627 ( .A0(n8057), .A1(n10609), .B0(n7367), .B1(n12120), .Y(n8053) );
  AOI22XLTS U5545 ( .A0(n10953), .A1(n6011), .B0(n10554), .B1(n5803), .Y(n6004) );
  AOI22XLTS U5312 ( .A0(n11711), .A1(n11970), .B0(n12247), .B1(n12271), .Y(
        n5555) );
  OAI22XLTS U5306 ( .A0(n5543), .A1(n11313), .B0(n5387), .B1(n10469), .Y(n5542) );
  OAI211XLTS U5542 ( .A0(n12210), .A1(n5291), .B0(n6008), .C0(n6009), .Y(n6007) );
  OAI22XLTS U2229 ( .A0(n1662), .A1(n10176), .B0(n11949), .B1(n12563), .Y(
        n2949) );
  AOI32XLTS U5980 ( .A0(n9538), .A1(n10878), .A2(n5917), .B0(n10585), .B1(
        n10879), .Y(n6521) );
  OAI22XLTS U3607 ( .A0(n10419), .A1(n10817), .B0(n11399), .B1(n12397), .Y(
        n4118) );
  AOI31XLTS U5977 ( .A0(n6107), .A1(n10100), .A2(n10170), .B0(n6255), .Y(n6519) );
  OAI22XLTS U2201 ( .A0(n2891), .A1(n11435), .B0(n10676), .B1(n2924), .Y(n2922) );
  OAI22XLTS U5490 ( .A0(n10513), .A1(n10923), .B0(n11217), .B1(n12426), .Y(
        n5918) );
  AOI22XLTS U7751 ( .A0(n11880), .A1(n11033), .B0(n11633), .B1(n10669), .Y(
        n8150) );
  OR2X2TS U4942 ( .A(n11703), .B(n11249), .Y(n4303) );
  AOI22XLTS U3441 ( .A0(n11720), .A1(n12051), .B0(n12236), .B1(n12213), .Y(
        n3800) );
  OAI22XLTS U5557 ( .A0(n10983), .A1(n9965), .B0(n10825), .B1(n10980), .Y(
        n6036) );
  OAI22XLTS U3435 ( .A0(n3788), .A1(n11292), .B0(n3589), .B1(n10437), .Y(n3787) );
  OAI22XLTS U2126 ( .A0(n2815), .A1(n11429), .B0(n10663), .B1(n2848), .Y(n2846) );
  AOI32XLTS U4097 ( .A0(n9451), .A1(n10889), .A2(n4117), .B0(n10408), .B1(
        n10888), .Y(n4721) );
  OAI211XLTS U7218 ( .A0(n7426), .A1(n10042), .B0(n7427), .C0(n7428), .Y(n7411) );
  AOI22XLTS U7917 ( .A0(n11914), .A1(n11516), .B0(n12349), .B1(n11123), .Y(
        n8320) );
  AOI31XLTS U7360 ( .A0(sa31[1]), .A1(n9869), .A2(n10077), .B0(n7728), .Y(
        n7722) );
  AOI22XLTS U7359 ( .A0(n11896), .A1(n11125), .B0(n9866), .B1(n11151), .Y(
        n7723) );
  INVX1TS U2047 ( .A(n2151), .Y(n2073) );
  OAI22XLTS U3643 ( .A0(n3550), .A1(n10911), .B0(n3868), .B1(n11243), .Y(n4175) );
  AOI32XLTS U2390 ( .A0(n11446), .A1(n3082), .A2(n10621), .B0(n10524), .B1(
        n3082), .Y(n3081) );
  OAI22XLTS U1971 ( .A0(n11584), .A1(n11149), .B0(n10982), .B1(n11435), .Y(
        n2700) );
  OAI22XLTS U2646 ( .A0(n11889), .A1(n10982), .B0(n12475), .B1(n1863), .Y(
        n3170) );
  AOI22XLTS U7873 ( .A0(n7313), .A1(n11927), .B0(n11592), .B1(n11140), .Y(
        n8279) );
  OAI22XLTS U3670 ( .A0(n9654), .A1(n10113), .B0(n10472), .B1(n4221), .Y(n4220) );
  INVX1TS U8447 ( .A(n7123), .Y(n8092) );
  OAI211XLTS U1804 ( .A0(n11859), .A1(n10960), .B0(n2481), .C0(n2482), .Y(
        n2479) );
  AOI22XLTS U5513 ( .A0(n6337), .A1(n5962), .B0(n10181), .B1(n5670), .Y(n5960)
         );
  OAI22XLTS U1958 ( .A0(n11478), .A1(n10275), .B0(n10208), .B1(n11899), .Y(
        n2681) );
  OAI22XLTS U1806 ( .A0(n11459), .A1(n10192), .B0(n10621), .B1(n10592), .Y(
        n2478) );
  OAI22XLTS U2882 ( .A0(n9109), .A1(n10215), .B0(n2431), .B1(n10255), .Y(n3248) );
  AOI32XLTS U7580 ( .A0(n9849), .A1(n11145), .A2(sa31[2]), .B0(n11098), .B1(
        n11144), .Y(n8010) );
  OAI22XLTS U1807 ( .A0(n11851), .A1(n10188), .B0(n11015), .B1(n11075), .Y(
        n2477) );
  OAI22XLTS U2807 ( .A0(n2844), .A1(n12469), .B0(n2805), .B1(n10993), .Y(n3216) );
  OAI22XLTS U3886 ( .A0(n12569), .A1(n11713), .B0(n10872), .B1(n12412), .Y(
        n4487) );
  OAI22XLTS U3671 ( .A0(n3589), .A1(n10893), .B0(n3893), .B1(n11238), .Y(n4219) );
  OAI22XLTS U3723 ( .A0(n11762), .A1(n12023), .B0(n10871), .B1(n10792), .Y(
        n4295) );
  CLKINVX2TS U4401 ( .A(n4021), .Y(n3837) );
  OAI22XLTS U5667 ( .A0(n10820), .A1(n11673), .B0(n12209), .B1(n10186), .Y(
        n6178) );
  AND2X2TS U2634 ( .A(n11900), .B(n12353), .Y(n1728) );
  INVX1TS U7928 ( .A(n7828), .Y(n7485) );
  OAI22XLTS U5590 ( .A0(n9714), .A1(n10210), .B0(n10427), .B1(n6087), .Y(n6086) );
  OAI22XLTS U7532 ( .A0(n11467), .A1(n10664), .B0(n11540), .B1(n11830), .Y(
        n7948) );
  OAI31XLTS U5646 ( .A0(n10416), .A1(n6049), .A2(n9986), .B0(n6160), .Y(n6159)
         );
  OAI22XLTS U1972 ( .A0(n11625), .A1(n10267), .B0(n11901), .B1(n11483), .Y(
        n2699) );
  CLKBUFX2TS U4251 ( .A(n12569), .Y(n3917) );
  OAI22XLTS U3642 ( .A0(n9658), .A1(n10106), .B0(n10490), .B1(n4177), .Y(n4176) );
  OAI22XLTS U5591 ( .A0(n5348), .A1(n5440), .B0(n5698), .B1(n11385), .Y(n6085)
         );
  OAI22XLTS U1973 ( .A0(n1725), .A1(n12176), .B0(n11899), .B1(n11436), .Y(
        n2698) );
  OAI22XLTS U5510 ( .A0(n11018), .A1(n11982), .B0(n12004), .B1(n10226), .Y(
        n5952) );
  OR2X2TS U8499 ( .A(n11535), .B(n10321), .Y(n7359) );
  NAND2XLTS U6464 ( .A(n10529), .B(n10428), .Y(n6089) );
  CLKBUFX2TS U8162 ( .A(n12617), .Y(n7698) );
  OAI22XLTS U2843 ( .A0(n11865), .A1(n10997), .B0(n12459), .B1(n12086), .Y(
        n3230) );
  OAI22XLTS U2685 ( .A0(n9112), .A1(n10207), .B0(n2387), .B1(n10279), .Y(n3188) );
  OAI22XLTS U2015 ( .A0(n1763), .A1(n12166), .B0(n11875), .B1(n11430), .Y(
        n2731) );
  AOI31XLTS U7324 ( .A0(n9850), .A1(n12183), .A2(n9854), .B0(n7657), .Y(n7640)
         );
  OAI22XLTS U2014 ( .A0(n11606), .A1(n10243), .B0(n11877), .B1(n11472), .Y(
        n2732) );
  OAI22XLTS U5618 ( .A0(n9718), .A1(n10218), .B0(n10444), .B1(n6131), .Y(n6130) );
  AND2X2TS U2831 ( .A(n11876), .B(n12348), .Y(n1766) );
  OAI22XLTS U5619 ( .A0(n5387), .A1(n5506), .B0(n5723), .B1(n11390), .Y(n6129)
         );
  CLKINVX2TS U6282 ( .A(n5807), .Y(n5632) );
  AOI21XLTS U1651 ( .A0(n11949), .A1(n11046), .B0(n10287), .Y(n2209) );
  AOI22XLTS U1997 ( .A0(n11117), .A1(n1933), .B0(n11929), .B1(n11566), .Y(
        n2718) );
  OAI31XLTS U3763 ( .A0(n10498), .A1(n4282), .A2(n9926), .B0(n4357), .Y(n4356)
         );
  OAI22XLTS U3890 ( .A0(n12568), .A1(n9640), .B0(n10782), .B1(n11774), .Y(
        n4499) );
  AOI31XLTS U8644 ( .A0(n10001), .A1(n10040), .A2(n11635), .B0(n7088), .Y(
        n8637) );
  OAI22XLTS U2000 ( .A0(n11466), .A1(n10251), .B0(n10216), .B1(n11875), .Y(
        n2714) );
  OAI22XLTS U2013 ( .A0(n11572), .A1(n11127), .B0(n10998), .B1(n11429), .Y(
        n2733) );
  AOI22XLTS U1955 ( .A0(n11137), .A1(n1870), .B0(n11942), .B1(n11578), .Y(
        n2685) );
  OAI22XLTS U1652 ( .A0(n10007), .A1(n12160), .B0(n12563), .B1(n11588), .Y(
        n2208) );
  OAI211XLTS U3837 ( .A0(n4099), .A1(n10821), .B0(n4436), .C0(n4437), .Y(n4435) );
  OAI21XLTS U7971 ( .A0(n10086), .A1(n11177), .B0(n8363), .Y(n8362) );
  OR2X2TS U8512 ( .A(n11160), .B(n8047), .Y(n7121) );
  OAI211XLTS U5478 ( .A0(n10874), .A1(n11365), .B0(n5897), .C0(n5898), .Y(
        n5891) );
  OAI31XLTS U5820 ( .A0(n6373), .A1(sa01[3]), .A2(n11990), .B0(n6294), .Y(
        n6361) );
  OAI22XLTS U4865 ( .A0(n4578), .A1(n12569), .B0(n3967), .B1(n12541), .Y(n5063) );
  OAI22XLTS U7551 ( .A0(n12158), .A1(n12128), .B0(n11574), .B1(n10085), .Y(
        n7968) );
  CLKINVX2TS U2337 ( .A(n1961), .Y(n2781) );
  OAI31XLTS U5744 ( .A0(n6265), .A1(n5366), .A2(n10469), .B0(n6266), .Y(n6260)
         );
  OAI22XLTS U2046 ( .A0(n2153), .A1(n10191), .B0(n2073), .B1(n11034), .Y(n2763) );
  NOR3XLTS U5945 ( .A(n9420), .B(n9424), .C(n10930), .Y(n6485) );
  OAI211XLTS U7552 ( .A0(n11166), .A1(n11118), .B0(n7971), .C0(n7289), .Y(
        n7961) );
  AOI32XLTS U2451 ( .A0(n9931), .A1(n3118), .A2(n10607), .B0(n10954), .B1(
        n3118), .Y(n3117) );
  OAI22XLTS U3633 ( .A0(n4160), .A1(n12008), .B0(n3866), .B1(n10844), .Y(n4156) );
  AOI21XLTS U3725 ( .A0(n10770), .A1(n10861), .B0(n11756), .Y(n4293) );
  OAI22XLTS U5947 ( .A0(n10929), .A1(n10452), .B0(n10918), .B1(n9774), .Y(
        n6493) );
  AOI32XLTS U8706 ( .A0(n11468), .A1(n8129), .A2(n10294), .B0(n12150), .B1(
        n8129), .Y(n8663) );
  AOI31XLTS U4432 ( .A0(n10882), .A1(n10368), .A2(n4281), .B0(n4732), .Y(n4934) );
  OAI211XLTS U3741 ( .A0(n11775), .A1(n10769), .B0(n4331), .C0(n4332), .Y(
        n4330) );
  OAI31XLTS U6616 ( .A0(sa23[1]), .A1(n9448), .A2(n9775), .B0(n5556), .Y(n6828) );
  OAI211XLTS U3801 ( .A0(n4043), .A1(n10848), .B0(n4396), .C0(n4397), .Y(n4395) );
  OAI211XLTS U2269 ( .A0(n11046), .A1(n9932), .B0(n2983), .C0(n2008), .Y(n2982) );
  AOI31XLTS U7827 ( .A0(n9894), .A1(n11180), .A2(n7594), .B0(n8177), .Y(n8236)
         );
  OAI22XLTS U7831 ( .A0(n7585), .A1(n11653), .B0(n11176), .B1(n12163), .Y(
        n8232) );
  OAI211XLTS U6121 ( .A0(n11735), .A1(n11992), .B0(n6647), .C0(n6648), .Y(
        n6646) );
  AOI211XLTS U8008 ( .A0(n12635), .A1(n7296), .B0(n8396), .C0(n8397), .Y(n8394) );
  AOI31XLTS U5806 ( .A0(sa01[1]), .A1(n9738), .A2(n10546), .B0(n6350), .Y(
        n6343) );
  OAI22XLTS U3885 ( .A0(n3910), .A1(n4807), .B0(n10111), .B1(n12024), .Y(n4488) );
  INVX1TS U5309 ( .A(n5523), .Y(n5546) );
  NAND3XLTS U2484 ( .A(n10606), .B(n12564), .C(n10695), .Y(n3126) );
  AOI31XLTS U4386 ( .A0(n10502), .A1(n12037), .A2(n10921), .B0(n10943), .Y(
        n4930) );
  OAI211XLTS U6085 ( .A0(n12019), .A1(n11729), .B0(n5652), .C0(n6612), .Y(
        n6608) );
  NOR2XLTS U3733 ( .A(n4319), .B(n12533), .Y(n4316) );
  OAI211XLTS U4270 ( .A0(n4503), .A1(n12382), .B0(n4874), .C0(n4875), .Y(n4873) );
  AOI22XLTS U1786 ( .A0(n11494), .A1(n1935), .B0(n11095), .B1(n9058), .Y(n2451) );
  OAI21XLTS U3700 ( .A0(n4261), .A1(n10754), .B0(n4262), .Y(n4250) );
  NOR2XLTS U2240 ( .A(n9959), .B(n11642), .Y(n2954) );
  AND2X2TS U7996 ( .A(n10046), .B(n12129), .Y(n7459) );
  OAI211XLTS U3389 ( .A0(n9901), .A1(n11380), .B0(n3660), .C0(n3661), .Y(n3657) );
  OAI22XLTS U4493 ( .A0(n4064), .A1(n12404), .B0(n4584), .B1(n10843), .Y(n4953) );
  OAI211XLTS U1516 ( .A0(n11882), .A1(n11877), .B0(n1902), .C0(n1903), .Y(
        n1899) );
  OAI211XLTS U3562 ( .A0(n3685), .A1(n11260), .B0(n4041), .C0(n4042), .Y(n4035) );
  OR2X2TS U8472 ( .A(n11443), .B(n10017), .Y(n7364) );
  OAI22XLTS U4490 ( .A0(n4595), .A1(n11244), .B0(n4161), .B1(n10109), .Y(n4954) );
  OAI22XLTS U5258 ( .A0(n5413), .A1(n12494), .B0(n5414), .B1(n10153), .Y(n5408) );
  AOI31XLTS U7224 ( .A0(n9505), .A1(n10273), .A2(n7440), .B0(n7441), .Y(n7433)
         );
  OAI22XLTS U2444 ( .A0(n2533), .A1(n11589), .B0(n10690), .B1(n11643), .Y(
        n3112) );
  OAI22XLTS U3002 ( .A0(n2465), .A1(n11034), .B0(n2769), .B1(n11448), .Y(n3273) );
  OAI22XLTS U4473 ( .A0(n4160), .A1(n10839), .B0(n11411), .B1(n11344), .Y(
        n4947) );
  AOI31XLTS U3387 ( .A0(n9678), .A1(n9674), .A2(n12411), .B0(n10859), .Y(n3645) );
  AOI32XLTS U1879 ( .A0(n2586), .A1(n10615), .A2(n9844), .B0(n11005), .B1(
        n10616), .Y(n2585) );
  OAI31XLTS U3826 ( .A0(n4422), .A1(n3529), .A2(n10446), .B0(n4423), .Y(n4417)
         );
  OAI22XLTS U3989 ( .A0(n10837), .A1(n10482), .B0(n10848), .B1(n9668), .Y(
        n4621) );
  INVX1TS U7926 ( .A(n7681), .Y(n7330) );
  OAI211XLTS U5683 ( .A0(n5843), .A1(n10890), .B0(n6199), .C0(n6200), .Y(n6198) );
  AOI22XLTS U3917 ( .A0(n11374), .A1(n4325), .B0(n10460), .B1(n4536), .Y(n4535) );
  OAI22XLTS U2805 ( .A0(n9108), .A1(n11429), .B0(n2246), .B1(n10992), .Y(n3217) );
  OAI22XLTS U3635 ( .A0(n4161), .A1(n11339), .B0(n9915), .B1(n10839), .Y(n4154) );
  AOI22XLTS U7657 ( .A0(n10320), .A1(n12089), .B0(n11628), .B1(n12312), .Y(
        n8077) );
  CLKINVX1TS U8001 ( .A(n8179), .Y(n8370) );
  INVX1TS U8315 ( .A(n7963), .Y(n8529) );
  AOI31XLTS U1630 ( .A0(n10360), .A1(n2167), .A2(n10588), .B0(n2169), .Y(n2156) );
  OAI211XLTS U7800 ( .A0(n10049), .A1(n11183), .B0(n8200), .C0(n8201), .Y(
        n8199) );
  CLKINVX2TS U2892 ( .A(n1935), .Y(n2272) );
  NAND4XLTS U4205 ( .A(n4814), .B(n4815), .C(n4485), .D(n4291), .Y(n4809) );
  AOI31XLTS U8757 ( .A0(n9624), .A1(sa20[2]), .A2(n10274), .B0(n8114), .Y(
        n8677) );
  OAI22XLTS U6104 ( .A0(n6631), .A1(n12011), .B0(n6632), .B1(n10234), .Y(n6628) );
  OAI22XLTS U3376 ( .A0(n3615), .A1(n12546), .B0(n3616), .B1(n9907), .Y(n3610)
         );
  OAI211XLTS U4199 ( .A0(n12412), .A1(n9641), .B0(n4812), .C0(n3922), .Y(n4811) );
  OAI22XLTS U7717 ( .A0(n7069), .A1(n10297), .B0(n11819), .B1(n9467), .Y(n8125) );
  INVX1TS U7780 ( .A(n8123), .Y(n8162) );
  OAI211XLTS U2273 ( .A0(n10689), .A1(n11949), .B0(n2985), .C0(n2610), .Y(
        n2981) );
  OAI211XLTS U3595 ( .A0(n10894), .A1(n11255), .B0(n4097), .C0(n4098), .Y(
        n4091) );
  OAI211XLTS U7916 ( .A0(n10647), .A1(n11902), .B0(n8320), .C0(n8321), .Y(
        n8319) );
  OAI21XLTS U2281 ( .A0(n9995), .A1(n12554), .B0(n2606), .Y(n2993) );
  INVX1TS U7841 ( .A(n8250), .Y(n8210) );
  OAI22XLTS U7711 ( .A0(n8123), .A1(n10594), .B0(n7216), .B1(n11838), .Y(n8119) );
  OAI22XLTS U7076 ( .A0(n7069), .A1(n11420), .B0(n7071), .B1(n11426), .Y(n7062) );
  OAI211XLTS U6774 ( .A0(n9723), .A1(n9710), .B0(n6672), .C0(n6881), .Y(n6880)
         );
  OAI22XLTS U5583 ( .A0(n6071), .A1(n11264), .B0(n9945), .B1(n10902), .Y(n6064) );
  OAI22XLTS U6748 ( .A0(n5958), .A1(n10976), .B0(n6378), .B1(n11748), .Y(n6861) );
  CLKINVX1TS U5669 ( .A(n6186), .Y(n6185) );
  AOI31XLTS U5340 ( .A0(n9816), .A1(n5625), .A2(n11341), .B0(n5627), .Y(n5624)
         );
  OAI22XLTS U8691 ( .A0(n8123), .A1(n11770), .B0(n11469), .B1(n8127), .Y(n8656) );
  AOI31XLTS U3606 ( .A0(n4117), .A1(n11986), .A2(n11191), .B0(n4118), .Y(n4114) );
  AOI31XLTS U5456 ( .A0(n5861), .A1(n12034), .A2(n11186), .B0(n5862), .Y(n5858) );
  OAI22XLTS U6373 ( .A0(n6395), .A1(n11385), .B0(n6071), .B1(n10213), .Y(n6753) );
  OAI22XLTS U5609 ( .A0(n6114), .A1(n12040), .B0(n5721), .B1(n10925), .Y(n6110) );
  INVX1TS U4346 ( .A(n4261), .Y(n4784) );
  OAI22XLTS U7594 ( .A0(n11903), .A1(n10342), .B0(n7829), .B1(n11108), .Y(
        n8028) );
  OAI22XLTS U6376 ( .A0(n5864), .A1(n12416), .B0(n10462), .B1(n10896), .Y(
        n6752) );
  OAI22XLTS U3661 ( .A0(n4204), .A1(n11993), .B0(n3891), .B1(n10817), .Y(n4200) );
  OAI31XLTS U4538 ( .A0(sa11[1]), .A1(n9244), .A2(n9669), .B0(n3735), .Y(n4971) );
  AOI31XLTS U7477 ( .A0(sa13[1]), .A1(n7550), .A2(n10262), .B0(n7881), .Y(
        n7875) );
  AOI22XLTS U1759 ( .A0(n11488), .A1(n1872), .B0(n11111), .B1(n9065), .Y(n2407) );
  OAI211XLTS U4916 ( .A0(n12567), .A1(n10770), .B0(n5097), .C0(n4559), .Y(
        n5096) );
  OAI22XLTS U4064 ( .A0(n10809), .A1(n10463), .B0(n10822), .B1(n9671), .Y(
        n4693) );
  OAI31XLTS U7590 ( .A0(n9370), .A1(n11101), .A2(n8022), .B0(n7643), .Y(n8021)
         );
  OAI31XLTS U6421 ( .A0(sa12[1]), .A1(n9440), .A2(n9771), .B0(n5490), .Y(n6770) );
  AOI21XLTS U3545 ( .A0(n10756), .A1(n10403), .B0(n11805), .Y(n4010) );
  AOI31XLTS U7598 ( .A0(n7835), .A1(n11523), .A2(n12356), .B0(n10707), .Y(
        n8019) );
  OAI22XLTS U7600 ( .A0(n7828), .A1(n10647), .B0(n7494), .B1(n11609), .Y(n8030) );
  AOI21XLTS U6027 ( .A0(n11979), .A1(n10834), .B0(n5637), .Y(n6563) );
  OR2X2TS U7354 ( .A(n11856), .B(n11551), .Y(n7335) );
  OAI31XLTS U6806 ( .A0(n10722), .A1(n11018), .A2(n6897), .B0(n6898), .Y(n6894) );
  NOR3XLTS U5870 ( .A(n9411), .B(n9415), .C(n10903), .Y(n6413) );
  AOI31XLTS U6314 ( .A0(n11228), .A1(n10327), .A2(n6738), .B0(n6532), .Y(n6733) );
  OAI31XLTS U5708 ( .A0(n6225), .A1(n5327), .A2(n10462), .B0(n6226), .Y(n6220)
         );
  OAI22XLTS U5581 ( .A0(n6070), .A1(n12026), .B0(n5696), .B1(n10898), .Y(n6066) );
  OAI211XLTS U7308 ( .A0(n12162), .A1(n11574), .B0(n7612), .C0(n7613), .Y(
        n7600) );
  OAI22XLTS U5893 ( .A0(n10530), .A1(n11204), .B0(n10902), .B1(n10857), .Y(
        n6441) );
  OAI22XLTS U4125 ( .A0(n4386), .A1(n12387), .B0(n3985), .B1(n10119), .Y(n4739) );
  AOI211XLTS U6036 ( .A0(n10840), .A1(n11980), .B0(n6572), .C0(n6573), .Y(
        n6567) );
  AOI31XLTS U6267 ( .A0(n10824), .A1(n11976), .A2(n10846), .B0(n10819), .Y(
        n6729) );
  OAI211XLTS U7403 ( .A0(n12328), .A1(n10594), .B0(n7785), .C0(n7050), .Y(
        n7781) );
  OAI211XLTS U7400 ( .A0(n12068), .A1(n10618), .B0(n7783), .C0(n7380), .Y(
        n7782) );
  OAI22XLTS U2194 ( .A0(n2313), .A1(n11476), .B0(n2891), .B1(n10212), .Y(n2916) );
  AOI31XLTS U1888 ( .A0(n2598), .A1(n1671), .A2(n2599), .B0(n2600), .Y(n2596)
         );
  INVX1TS U5284 ( .A(n5457), .Y(n5480) );
  OAI31XLTS U3862 ( .A0(n4462), .A1(n3568), .A2(n10438), .B0(n4463), .Y(n4457)
         );
  OAI211XLTS U5445 ( .A0(n10858), .A1(n11361), .B0(n5841), .C0(n5842), .Y(
        n5835) );
  OAI31XLTS U4733 ( .A0(sa22[1]), .A1(n9252), .A2(n9671), .B0(n3801), .Y(n5029) );
  INVX1TS U8633 ( .A(n7069), .Y(n8158) );
  AND2X2TS U1903 ( .A(n10607), .B(n9701), .Y(n1823) );
  CLKINVX2TS U2695 ( .A(n1872), .Y(n2339) );
  AOI21XLTS U5421 ( .A0(n10991), .A1(n10522), .B0(n11691), .Y(n5794) );
  AOI22XLTS U7911 ( .A0(n12634), .A1(n11862), .B0(n12189), .B1(n11591), .Y(
        n8312) );
  OAI22XLTS U6747 ( .A0(n6374), .A1(n11728), .B0(n5746), .B1(n9723), .Y(n6862)
         );
  AOI31XLTS U5489 ( .A0(n5917), .A1(n12049), .A2(sa23[2]), .B0(n5918), .Y(
        n5914) );
  AOI31XLTS U3458 ( .A0(sa33[2]), .A1(n3830), .A2(n11266), .B0(n3832), .Y(
        n3829) );
  INVX1TS U6228 ( .A(n6028), .Y(n6584) );
  OAI22XLTS U4085 ( .A0(n10382), .A1(n11399), .B0(n10809), .B1(n10893), .Y(
        n4713) );
  AOI211XLTS U8455 ( .A0(n10605), .A1(n10018), .B0(n8573), .C0(n7261), .Y(
        n8572) );
  AOI22XLTS U2173 ( .A0(n12599), .A1(n9064), .B0(n11105), .B1(n10552), .Y(
        n2897) );
  OAI22XLTS U4109 ( .A0(n12549), .A1(n10151), .B0(n11804), .B1(n9920), .Y(
        n4733) );
  AOI22XLTS U7583 ( .A0(n12189), .A1(n11896), .B0(n11860), .B1(n11150), .Y(
        n8007) );
  OAI22XLTS U3663 ( .A0(n4205), .A1(n11291), .B0(n9911), .B1(n10811), .Y(n4198) );
  NOR3XLTS U4062 ( .A(n9218), .B(n9221), .C(n10810), .Y(n4685) );
  AOI31XLTS U3573 ( .A0(n4061), .A1(n12003), .A2(sa11[2]), .B0(n4062), .Y(
        n4058) );
  OAI22XLTS U5872 ( .A0(n10902), .A1(n10435), .B0(n10890), .B1(n9770), .Y(
        n6421) );
  OAI21XLTS U4893 ( .A0(n12492), .A1(n10866), .B0(n5086), .Y(n5085) );
  OAI22XLTS U6356 ( .A0(n6070), .A1(n10904), .B0(n11205), .B1(n11257), .Y(
        n6746) );
  AOI22XLTS U1656 ( .A0(n10584), .A1(n2221), .B0(n11507), .B1(n2222), .Y(n2218) );
  CLKINVX1TS U3786 ( .A(n4382), .Y(n4381) );
  INVX1TS U6823 ( .A(n5759), .Y(n6335) );
  OAI22XLTS U5611 ( .A0(n6115), .A1(n11312), .B0(n9949), .B1(n10931), .Y(n6108) );
  OAI22XLTS U7094 ( .A0(n7123), .A1(n11802), .B0(n7125), .B1(n12081), .Y(n7116) );
  OAI21XLTS U5552 ( .A0(n6028), .A1(n10989), .B0(n6029), .Y(n6018) );
  OAI31XLTS U4919 ( .A0(n10318), .A1(n10790), .A2(n5098), .B0(n5099), .Y(n5095) );
  AOI21XLTS U4144 ( .A0(n11809), .A1(n10932), .B0(n3842), .Y(n4763) );
  OAI22XLTS U6750 ( .A0(n6632), .A1(n11984), .B0(n5763), .B1(n12287), .Y(n6860) );
  AOI32XLTS U6782 ( .A0(n11371), .A1(n6673), .A2(n11989), .B0(n10229), .B1(
        n6673), .Y(n6887) );
  INVX1TS U3438 ( .A(n3768), .Y(n3791) );
  NOR3XLTS U3987 ( .A(n9211), .B(n9214), .C(n10838), .Y(n4613) );
  CLKINVX2TS U4884 ( .A(n4536), .Y(n3913) );
  OAI31XLTS U6762 ( .A0(sa01[7]), .A1(n6872), .A2(n11372), .B0(n6873), .Y(
        n6871) );
  INVX1TS U3413 ( .A(n3702), .Y(n3725) );
  OAI22XLTS U5754 ( .A0(n12014), .A1(n5579), .B0(n6277), .B1(n11754), .Y(n6275) );
  OAI211XLTS U7910 ( .A0(n11611), .A1(n11902), .B0(n8312), .C0(n8313), .Y(
        n8311) );
  OAI22XLTS U1622 ( .A0(n10629), .A1(n10593), .B0(n11548), .B1(n11073), .Y(
        n2147) );
  OAI22XLTS U3958 ( .A0(n11350), .A1(n11260), .B0(n9135), .B1(n12446), .Y(
        n4585) );
  OAI211XLTS U4142 ( .A0(n10403), .A1(n12388), .B0(n4763), .C0(n4370), .Y(
        n4762) );
  OAI211XLTS U7410 ( .A0(n10041), .A1(n11843), .B0(n7794), .C0(n7795), .Y(
        n7793) );
  OAI211XLTS U8010 ( .A0(n11639), .A1(n11950), .B0(n8398), .C0(n8256), .Y(
        n8392) );
  OAI22XLTS U5839 ( .A0(n6068), .A1(n9946), .B0(n5694), .B1(n11383), .Y(n6387)
         );
  CLKINVX2TS U2401 ( .A(n2213), .Y(n1809) );
  OAI211XLTS U1996 ( .A0(n12168), .A1(n11607), .B0(n2717), .C0(n2718), .Y(
        n2716) );
  AOI2BB2XLTS U6414 ( .B0(n11211), .B1(n9298), .A0N(n11253), .A1N(n6068), .Y(
        n6772) );
  OAI31XLTS U2045 ( .A0(sa03[3]), .A1(n2765), .A2(n11079), .B0(n2766), .Y(
        n2764) );
  OAI211XLTS U8007 ( .A0(n12172), .A1(n11182), .B0(n8394), .C0(n8395), .Y(
        n8393) );
  NAND3XLTS U2293 ( .A(n3001), .B(n2559), .C(n3002), .Y(n2614) );
  OAI22XLTS U3912 ( .A0(n9641), .A1(n4480), .B0(n12381), .B1(n11755), .Y(n4530) );
  OAI211XLTS U7276 ( .A0(n10266), .A1(n12103), .B0(n7543), .C0(n7544), .Y(
        n7542) );
  OAI22XLTS U5841 ( .A0(n11251), .A1(n11361), .B0(n9330), .B1(n12386), .Y(
        n6385) );
  AOI31XLTS U5517 ( .A0(n12680), .A1(n9739), .A2(n9977), .B0(n5968), .Y(n5965)
         );
  OAI22XLTS U4150 ( .A0(n10120), .A1(n10108), .B0(n10402), .B1(n10938), .Y(
        n4771) );
  NAND2XLTS U3035 ( .A(n11440), .B(n11562), .Y(n3296) );
  AOI2BB2XLTS U6609 ( .B0(n11223), .B1(n9308), .A0N(n11300), .A1N(n6112), .Y(
        n6830) );
  OAI22XLTS U3956 ( .A0(n4158), .A1(n9916), .B0(n3864), .B1(n11242), .Y(n4587)
         );
  OAI211XLTS U7709 ( .A0(n7425), .A1(n12150), .B0(n8121), .C0(n8122), .Y(n8120) );
  OAI211XLTS U2153 ( .A0(n10543), .A1(n11618), .B0(n2878), .C0(n2879), .Y(
        n2877) );
  OAI211XLTS U7504 ( .A0(n12067), .A1(n11844), .B0(n7915), .C0(n7916), .Y(
        n7914) );
  OAI31XLTS U4588 ( .A0(n9358), .A1(n4422), .A2(n10447), .B0(n4077), .Y(n4991)
         );
  AOI31XLTS U2443 ( .A0(sa32[4]), .A1(n12152), .A2(n2560), .B0(n3112), .Y(
        n3110) );
  OAI22XLTS U5665 ( .A0(n5427), .A1(n9966), .B0(n10521), .B1(n10830), .Y(n6180) );
  AOI21XLTS U3386 ( .A0(n3647), .A1(n10871), .B0(n10865), .Y(n3646) );
  OAI211XLTS U2172 ( .A0(n2895), .A1(n11484), .B0(n2896), .C0(n2897), .Y(n2894) );
  AOI32XLTS U8434 ( .A0(n12122), .A1(n8557), .A2(n12558), .B0(n11873), .B1(
        n8557), .Y(n8552) );
  AOI31XLTS U3979 ( .A0(n10910), .A1(n11363), .A2(n3864), .B0(n11344), .Y(
        n4611) );
  OAI22XLTS U3724 ( .A0(n10144), .A1(n12538), .B0(n12208), .B1(n10455), .Y(
        n4294) );
  AOI31XLTS U5937 ( .A0(n10873), .A1(n11288), .A2(n5719), .B0(n11305), .Y(
        n6483) );
  OAI22XLTS U3529 ( .A0(n12282), .A1(n10108), .B0(n9914), .B1(n11805), .Y(
        n3983) );
  OAI211XLTS U8566 ( .A0(n10677), .A1(n12095), .B0(n8612), .C0(n7236), .Y(
        n8608) );
  OAI22XLTS U3660 ( .A0(n4202), .A1(n3595), .B0(n9161), .B1(n11297), .Y(n4201)
         );
  OAI22XLTS U7715 ( .A0(n7786), .A1(n10298), .B0(n7927), .B1(n10293), .Y(n8126) );
  AOI2BB2XLTS U4531 ( .B0(n11406), .B1(n9106), .A0N(n11352), .A1N(n4158), .Y(
        n4973) );
  OAI22XLTS U3782 ( .A0(n3629), .A1(n9914), .B0(n10402), .B1(n10938), .Y(n4376) );
  OAI22XLTS U5608 ( .A0(n6112), .A1(n5393), .B0(n9367), .B1(n11306), .Y(n6111)
         );
  CLKINVX2TS U8085 ( .A(n7491), .Y(n8306) );
  OAI211XLTS U7194 ( .A0(n11070), .A1(n11419), .B0(n7381), .C0(n7382), .Y(
        n7375) );
  OAI211XLTS U3882 ( .A0(n9674), .A1(n10777), .B0(n4490), .C0(n3966), .Y(n4489) );
  OAI211XLTS U2097 ( .A0(n2819), .A1(n11470), .B0(n2820), .C0(n2821), .Y(n2818) );
  OAI22XLTS U2987 ( .A0(n11446), .A1(n12098), .B0(n10510), .B1(n10625), .Y(
        n3266) );
  OAI22XLTS U7672 ( .A0(n7549), .A1(n11932), .B0(n7770), .B1(n12336), .Y(n8089) );
  OAI31XLTS U1878 ( .A0(n2558), .A1(n11637), .A2(n9044), .B0(n2585), .Y(n2578)
         );
  AOI32XLTS U5728 ( .A0(n11301), .A1(n6247), .A2(n10453), .B0(n10571), .B1(
        n6247), .Y(n6246) );
  OAI22XLTS U7405 ( .A0(n7786), .A1(n11842), .B0(n7787), .B1(n11425), .Y(n7780) );
  OAI211XLTS U2078 ( .A0(n10569), .A1(n11600), .B0(n2802), .C0(n2803), .Y(
        n2801) );
  OAI211XLTS U8752 ( .A0(n10293), .A1(n11777), .B0(n8677), .C0(n7164), .Y(
        n8673) );
  AOI22XLTS U7905 ( .A0(n11915), .A1(n7332), .B0(n11124), .B1(n7826), .Y(n8304) );
  OAI22XLTS U5580 ( .A0(n6068), .A1(n5354), .B0(n9359), .B1(n11259), .Y(n6067)
         );
  AOI31XLTS U4054 ( .A0(n10895), .A1(n11316), .A2(n3889), .B0(n11296), .Y(
        n4683) );
  OAI31XLTS U4878 ( .A0(n10319), .A1(n5074), .A2(n12207), .B0(n5075), .Y(n5073) );
  OAI31XLTS U2461 ( .A0(n2557), .A1(n12679), .A2(n1670), .B0(n3120), .Y(n3119)
         );
  OAI211XLTS U4240 ( .A0(n12532), .A1(n11775), .B0(n4848), .C0(n4849), .Y(
        n4847) );
  AOI2BB2XLTS U4726 ( .B0(n11394), .B1(n9115), .A0N(n11303), .A1N(n4202), .Y(
        n5031) );
  OAI211XLTS U2797 ( .A0(n12348), .A1(n12460), .B0(n3213), .C0(n2843), .Y(
        n3212) );
  OAI22XLTS U4031 ( .A0(n4202), .A1(n9912), .B0(n3889), .B1(n11236), .Y(n4659)
         );
  AOI32XLTS U3810 ( .A0(n11352), .A1(n4404), .A2(n10481), .B0(n10376), .B1(
        n4404), .Y(n4403) );
  NOR2XLTS U4899 ( .A(n10769), .B(n9670), .Y(n4566) );
  OAI31XLTS U7562 ( .A0(n7630), .A1(n9882), .A2(n10351), .B0(n7993), .Y(n7990)
         );
  AOI31XLTS U2392 ( .A0(n11015), .A1(n10509), .A2(n9923), .B0(n10593), .Y(
        n3080) );
  OAI211XLTS U1758 ( .A0(n2405), .A1(n12079), .B0(n2406), .C0(n2407), .Y(n2404) );
  OAI22XLTS U3754 ( .A0(n10163), .A1(n10765), .B0(n10945), .B1(n10107), .Y(
        n4347) );
  OAI211XLTS U1785 ( .A0(n2449), .A1(n12086), .B0(n2450), .C0(n2451), .Y(n2448) );
  OAI211XLTS U7793 ( .A0(n10745), .A1(n12164), .B0(n8188), .C0(n8189), .Y(
        n8186) );
  INVX1TS U7649 ( .A(n7766), .Y(n7513) );
  OAI22XLTS U3091 ( .A0(n10236), .A1(n11073), .B0(n11548), .B1(n12098), .Y(
        n3289) );
  OAI22XLTS U5637 ( .A0(n10412), .A1(n5630), .B0(n10820), .B1(n10205), .Y(
        n6150) );
  OAI22XLTS U5419 ( .A0(n10417), .A1(n10205), .B0(n12203), .B1(n10826), .Y(
        n5796) );
  OAI31XLTS U6471 ( .A0(sa12[7]), .A1(n6225), .A2(n10461), .B0(n5877), .Y(
        n6790) );
  OAI211XLTS U7625 ( .A0(n7535), .A1(n12335), .B0(n8055), .C0(n8056), .Y(n8054) );
  OAI211XLTS U2600 ( .A0(n12354), .A1(n12477), .B0(n3153), .C0(n2919), .Y(
        n3152) );
  OAI22XLTS U3632 ( .A0(n4158), .A1(n10482), .B0(n9154), .B1(n11346), .Y(n4157) );
  AND2X2TS U3026 ( .A(n11080), .B(n11458), .Y(n2057) );
  OAI22XLTS U6033 ( .A0(n10190), .A1(n10205), .B0(n10521), .B1(n10829), .Y(
        n6571) );
  AOI22XLTS U1650 ( .A0(n12187), .A1(n11953), .B0(n12093), .B1(n12182), .Y(
        n2211) );
  OAI211XLTS U8057 ( .A0(n11511), .A1(n10062), .B0(n8285), .C0(n8438), .Y(
        n8437) );
  OAI22XLTS U3543 ( .A0(n10499), .A1(n10107), .B0(n12282), .B1(n10504), .Y(
        n4012) );
  OAI22XLTS U5916 ( .A0(n11299), .A1(n11365), .B0(n9346), .B1(n12402), .Y(
        n6457) );
  AOI32XLTS U3846 ( .A0(n11304), .A1(n4444), .A2(n10464), .B0(n10371), .B1(
        n4444), .Y(n4443) );
  OAI31XLTS U4783 ( .A0(n9458), .A1(n4462), .A2(n10437), .B0(n4133), .Y(n5049)
         );
  OAI22XLTS U5914 ( .A0(n6112), .A1(n9950), .B0(n5719), .B1(n11389), .Y(n6459)
         );
  OAI211XLTS U6025 ( .A0(n10521), .A1(n12440), .B0(n6563), .C0(n6174), .Y(
        n6562) );
  OAI211XLTS U7203 ( .A0(n9802), .A1(n11794), .B0(n7401), .C0(n7402), .Y(n7400) );
  AOI211XLTS U4084 ( .A0(n4466), .A1(n10900), .B0(n4453), .C0(n4713), .Y(n4710) );
  AOI211XLTS U5892 ( .A0(n6229), .A1(n10852), .B0(n6216), .C0(n6441), .Y(n6438) );
  OAI31XLTS U6666 ( .A0(n9545), .A1(n6265), .A2(n10470), .B0(n5933), .Y(n6848)
         );
  INVX1TS U8657 ( .A(n7786), .Y(n7214) );
  AOI31XLTS U5862 ( .A0(n10857), .A1(n11239), .A2(n5694), .B0(n11257), .Y(
        n6411) );
  OAI31XLTS U1628 ( .A0(n10091), .A1(n9951), .A2(n11530), .B0(n2165), .Y(n2161) );
  OAI31XLTS U1817 ( .A0(n9855), .A1(n10960), .A2(n2508), .B0(n2509), .Y(n2506)
         );
  AOI211XLTS U1621 ( .A0(n12613), .A1(n11828), .B0(n2146), .C0(n2147), .Y(
        n2142) );
  AOI31XLTS U7719 ( .A0(n9813), .A1(n12149), .A2(n8127), .B0(n11419), .Y(n8124) );
  OAI211XLTS U4107 ( .A0(n12039), .A1(n10756), .B0(n3979), .C0(n4016), .Y(
        n4730) );
  OAI22XLTS U4862 ( .A0(n9938), .A1(n12573), .B0(n3962), .B1(n10455), .Y(n5065) );
  OAI31XLTS U6893 ( .A0(sa01[2]), .A1(n6351), .A2(n12285), .B0(n5945), .Y(
        n6856) );
  AOI31XLTS U2425 ( .A0(n10602), .A1(n12160), .A2(n1672), .B0(n10288), .Y(
        n3098) );
  NAND2XLTS U6787 ( .A(n10968), .B(n12299), .Y(n6889) );
  OAI211XLTS U4890 ( .A0(n10454), .A1(n10407), .B0(n4312), .C0(n4875), .Y(
        n5084) );
  OAI22XLTS U7223 ( .A0(n7065), .A1(n9501), .B0(n9798), .B1(n10594), .Y(n7437)
         );
  OAI22XLTS U3005 ( .A0(n3043), .A1(n10593), .B0(n2149), .B1(n11852), .Y(n3272) );
  OAI222XLTS U7246 ( .A0(n11902), .A1(n10660), .B0(n11521), .B1(n7489), .C0(
        n11510), .C1(n10651), .Y(n7481) );
  OAI22XLTS U2999 ( .A0(n2636), .A1(n12315), .B0(n2140), .B1(n11075), .Y(n3275) );
  AOI31XLTS U7635 ( .A0(n9826), .A1(n12335), .A2(n8061), .B0(n11800), .Y(n8058) );
  OAI211XLTS U4912 ( .A0(n4856), .A1(n12568), .B0(n5093), .C0(n4865), .Y(n3902) );
  AOI22XLTS U5799 ( .A0(n5574), .A1(n5974), .B0(n10478), .B1(n9407), .Y(n6339)
         );
  CLKINVX2TS U3085 ( .A(n3297), .Y(n2499) );
  OAI22XLTS U2362 ( .A0(n2750), .A1(n12099), .B0(n1964), .B1(n11447), .Y(n3057) );
  OAI31XLTS U7362 ( .A0(n10651), .A1(n7730), .A2(n7731), .B0(n7732), .Y(n7719)
         );
  CLKINVX2TS U1914 ( .A(n2630), .Y(n2060) );
  OAI211XLTS U1649 ( .A0(n9995), .A1(n11637), .B0(n2211), .C0(n2212), .Y(n2210) );
  OAI31XLTS U4341 ( .A0(n9888), .A1(n3507), .A2(n9657), .B0(n4911), .Y(n4908)
         );
  OAI211XLTS U8286 ( .A0(n8503), .A1(n10749), .B0(n8518), .C0(n8519), .Y(n8517) );
  NAND3XLTS U3899 ( .A(n10319), .B(n10115), .C(n4517), .Y(n4504) );
  AOI31XLTS U7561 ( .A0(n9565), .A1(sa02[1]), .A2(n10740), .B0(n7990), .Y(
        n7982) );
  OAI211XLTS U3571 ( .A0(n10398), .A1(n12445), .B0(n4058), .C0(n4059), .Y(
        n4056) );
  OAI31XLTS U1570 ( .A0(n2035), .A1(n2036), .A2(n10291), .B0(n2037), .Y(n2026)
         );
  OAI22XLTS U8069 ( .A0(n7850), .A1(n10651), .B0(n11522), .B1(n11866), .Y(
        n8444) );
  INVX1TS U3131 ( .A(n2750), .Y(n2159) );
  OAI22XLTS U7573 ( .A0(n11101), .A1(n9551), .B0(n11921), .B1(n11866), .Y(
        n8003) );
  OAI22XLTS U7608 ( .A0(n7659), .A1(n10074), .B0(n7833), .B1(n9858), .Y(n8035)
         );
  OAI31XLTS U6223 ( .A0(n9812), .A1(n5305), .A2(n9747), .B0(n6710), .Y(n6707)
         );
  OAI211XLTS U3604 ( .A0(n10389), .A1(n12427), .B0(n4114), .C0(n4115), .Y(
        n4112) );
  OAI211XLTS U5555 ( .A0(n10819), .A1(n6050), .B0(n6034), .C0(n6035), .Y(n6033) );
  OAI211XLTS U5487 ( .A0(n10536), .A1(n12401), .B0(n5914), .C0(n5915), .Y(
        n5912) );
  OAI211XLTS U8484 ( .A0(n11873), .A1(n9837), .B0(n7771), .C0(n8056), .Y(n8563) );
  CLKINVX2TS U3789 ( .A(n4348), .Y(n3628) );
  OAI211XLTS U1838 ( .A0(n9963), .A1(n1686), .B0(n1683), .C0(n2538), .Y(n2537)
         );
  OAI22XLTS U8478 ( .A0(n9825), .A1(n12115), .B0(n7246), .B1(n11848), .Y(n8581) );
  OAI2BB1XLTS U2292 ( .A0N(n2535), .A1N(n3000), .B0(n2614), .Y(n2999) );
  OAI22XLTS U2058 ( .A0(n2636), .A1(n11035), .B0(n2776), .B1(n11074), .Y(n2773) );
  OAI211XLTS U7904 ( .A0(n10723), .A1(n10660), .B0(n8304), .C0(n8305), .Y(
        n8303) );
  OAI211XLTS U5454 ( .A0(n5479), .A1(n12384), .B0(n5858), .C0(n5859), .Y(n5856) );
  OAI211XLTS U7547 ( .A0(n7963), .A1(n11950), .B0(n7965), .C0(n7966), .Y(n7962) );
  OAI211XLTS U2441 ( .A0(n3089), .A1(n10291), .B0(n3110), .C0(n2951), .Y(n3109) );
  OAI22XLTS U8663 ( .A0(n9814), .A1(n11818), .B0(n7174), .B1(n11831), .Y(n8645) );
  OAI31XLTS U1568 ( .A0(n9097), .A1(n9732), .A2(n9964), .B0(n2031), .Y(n2027)
         );
  OAI211XLTS U5623 ( .A0(n6134), .A1(n10537), .B0(n6135), .C0(n6136), .Y(n6123) );
  OAI22XLTS U4863 ( .A0(n4573), .A1(n12414), .B0(n3963), .B1(n10782), .Y(n5064) );
  OAI211XLTS U3655 ( .A0(n11314), .A1(n11994), .B0(n4194), .C0(n3577), .Y(
        n4193) );
  OAI211XLTS U6409 ( .A0(n10209), .A1(n10435), .B0(n6772), .C0(n6773), .Y(
        n6771) );
  OAI211XLTS U3558 ( .A0(n10849), .A1(n11346), .B0(n4037), .C0(n4038), .Y(
        n4036) );
  OAI211XLTS U5512 ( .A0(n5958), .A1(n10230), .B0(n5960), .C0(n5961), .Y(n5957) );
  OAI31XLTS U4165 ( .A0(sa33[1]), .A1(n9913), .A2(n4783), .B0(n3510), .Y(n4782) );
  OAI211XLTS U2150 ( .A0(n11631), .A1(n11901), .B0(n1860), .C0(n2873), .Y(
        n2872) );
  OAI211XLTS U3647 ( .A0(n4180), .A1(n3724), .B0(n4181), .C0(n4182), .Y(n4169)
         );
  AOI22XLTS U8049 ( .A0(n11957), .A1(n10729), .B0(n12191), .B1(n7712), .Y(
        n8433) );
  OAI211XLTS U5855 ( .A0(n10506), .A1(n12384), .B0(n6404), .C0(n5322), .Y(
        n6400) );
  NAND4XLTS U4471 ( .A(n4943), .B(n3852), .C(n4944), .D(n4945), .Y(n4942) );
  OAI211XLTS U2075 ( .A0(n11613), .A1(n11877), .B0(n1923), .C0(n2797), .Y(
        n2796) );
  NAND4XLTS U6354 ( .A(n6742), .B(n5682), .C(n6743), .D(n6744), .Y(n6741) );
  OAI211XLTS U2060 ( .A0(n2777), .A1(n10235), .B0(n1952), .C0(n2778), .Y(n2740) );
  AOI22XLTS U7077 ( .A0(n11431), .A1(n7074), .B0(n11031), .B1(n12457), .Y(
        n7061) );
  OAI22XLTS U5412 ( .A0(n5414), .A1(n10979), .B0(n5416), .B1(n10186), .Y(n5781) );
  OAI31XLTS U6124 ( .A0(n9824), .A1(n5589), .A2(n9397), .B0(n6650), .Y(n6645)
         );
  OAI211XLTS U5595 ( .A0(n6090), .A1(n10525), .B0(n6091), .C0(n6092), .Y(n6079) );
  NAND4XLTS U5909 ( .A(n5370), .B(n6452), .C(n6453), .D(n6454), .Y(n6451) );
  OAI211XLTS U4721 ( .A0(n10114), .A1(n10463), .B0(n5031), .C0(n5032), .Y(
        n5030) );
  OAI211XLTS U3627 ( .A0(n11362), .A1(n12009), .B0(n4150), .C0(n3538), .Y(
        n4149) );
  OAI22XLTS U7631 ( .A0(n9829), .A1(n11129), .B0(n7880), .B1(n10677), .Y(n8060) );
  OAI211XLTS U4755 ( .A0(n9110), .A1(n11290), .B0(n4210), .C0(n4225), .Y(n5039) );
  OAI31XLTS U2663 ( .A0(n9362), .A1(n3177), .A2(n10544), .B0(n3178), .Y(n3169)
         );
  OAI31XLTS U4243 ( .A0(n12671), .A1(n3639), .A2(n9683), .B0(n4851), .Y(n4846)
         );
  OAI22XLTS U6745 ( .A0(n5973), .A1(n12020), .B0(n5769), .B1(n10473), .Y(n6863) );
  AOI211XLTS U8477 ( .A0(n11445), .A1(n8065), .B0(n7743), .C0(n8581), .Y(n8565) );
  OAI22XLTS U5515 ( .A0(n5674), .A1(n11754), .B0(n5676), .B1(n10517), .Y(n5956) );
  NAND4XLTS U4026 ( .A(n3572), .B(n4652), .C(n4653), .D(n4654), .Y(n4651) );
  AOI31XLTS U8068 ( .A0(n10336), .A1(n8443), .A2(n12616), .B0(n8444), .Y(n8442) );
  OAI211XLTS U6638 ( .A0(n9302), .A1(n11312), .B0(n6120), .C0(n6135), .Y(n6838) );
  OAI211XLTS U1522 ( .A0(n11573), .A1(n10251), .B0(n1923), .C0(n1924), .Y(
        n1920) );
  AOI211XLTS U8662 ( .A0(n11033), .A1(n8131), .B0(n7774), .C0(n8645), .Y(n8642) );
  NAND4XLTS U1943 ( .A(n2081), .B(n2395), .C(n2675), .D(n2676), .Y(n2674) );
  OAI211XLTS U4047 ( .A0(n10419), .A1(n12428), .B0(n4676), .C0(n3563), .Y(
        n4672) );
  OAI211XLTS U5441 ( .A0(n10891), .A1(n11259), .B0(n5837), .C0(n5838), .Y(
        n5836) );
  OAI31XLTS U2860 ( .A0(n9282), .A1(n3237), .A2(n10570), .B0(n3238), .Y(n3229)
         );
  OAI211XLTS U1681 ( .A0(n12346), .A1(n10220), .B0(n2266), .C0(n2267), .Y(
        n2265) );
  OAI31XLTS U4925 ( .A0(n12671), .A1(n5102), .A2(n9675), .B0(n3641), .Y(n5100)
         );
  OAI22XLTS U5795 ( .A0(n5769), .A1(n10229), .B0(n5597), .B1(n6334), .Y(n6331)
         );
  OAI211XLTS U1441 ( .A0(n10676), .A1(n11632), .B0(n1704), .C0(n1705), .Y(
        n1701) );
  OAI211XLTS U1454 ( .A0(n10663), .A1(n11614), .B0(n1742), .C0(n1743), .Y(
        n1739) );
  OAI211XLTS U5526 ( .A0(n12014), .A1(n11728), .B0(n5985), .C0(n5986), .Y(
        n5980) );
  OAI211XLTS U5575 ( .A0(n11240), .A1(n12027), .B0(n6060), .C0(n5336), .Y(
        n6059) );
  OAI211XLTS U1620 ( .A0(n2140), .A1(n11834), .B0(n2142), .C0(n2143), .Y(n2139) );
  AOI211XLTS U7323 ( .A0(n12362), .A1(n12350), .B0(n7652), .C0(n7653), .Y(
        n7641) );
  OAI211XLTS U3457 ( .A0(n12387), .A1(n12066), .B0(n3828), .C0(n3829), .Y(
        n3826) );
  OAI211XLTS U1716 ( .A0(n12354), .A1(n10211), .B0(n2333), .C0(n2334), .Y(
        n2332) );
  NOR3XLTS U3732 ( .A(n4316), .B(n4317), .C(n4318), .Y(n4315) );
  NAND4XLTS U2785 ( .A(n3204), .B(n2106), .C(n2437), .D(n3205), .Y(n3203) );
  OAI22XLTS U3943 ( .A0(n3963), .A1(n10872), .B0(n4304), .B1(n10775), .Y(n4577) );
  CLKINVX1TS U1814 ( .A(n2502), .Y(n2500) );
  OAI22XLTS U3788 ( .A0(n3628), .A1(n10119), .B0(n3844), .B1(n10498), .Y(n4385) );
  OAI22XLTS U3913 ( .A0(n3963), .A1(n12491), .B0(n3647), .B1(n9677), .Y(n4529)
         );
  INVX1TS U3790 ( .A(n3987), .Y(n4384) );
  NAND4XLTS U5834 ( .A(n5331), .B(n6380), .C(n6381), .D(n6382), .Y(n6379) );
  NAND4XLTS U3951 ( .A(n3533), .B(n4580), .C(n4581), .D(n4582), .Y(n4579) );
  OAI22XLTS U7093 ( .A0(n7119), .A1(n10005), .B0(n9806), .B1(n12462), .Y(n7117) );
  OAI22XLTS U7268 ( .A0(n7119), .A1(n10053), .B0(n9806), .B1(n10608), .Y(n7525) );
  OAI211XLTS U7090 ( .A0(n12305), .A1(n12075), .B0(n7111), .C0(n7112), .Y(
        n7108) );
  OAI211XLTS U8614 ( .A0(n9814), .A1(n11772), .B0(n7930), .C0(n8617), .Y(n8616) );
  OAI211XLTS U4526 ( .A0(n10106), .A1(n10480), .B0(n4973), .C0(n4974), .Y(
        n4972) );
  OAI211XLTS U7072 ( .A0(n12067), .A1(n11765), .B0(n7057), .C0(n7058), .Y(
        n7054) );
  OAI31XLTS U6815 ( .A0(n10225), .A1(sa01[1]), .A2(n6900), .B0(n5591), .Y(
        n6899) );
  OAI22XLTS U2244 ( .A0(n2534), .A1(n9967), .B0(n2014), .B1(n11644), .Y(n2959)
         );
  OAI211XLTS U5339 ( .A0(n12439), .A1(n12196), .B0(n5623), .C0(n5624), .Y(
        n5621) );
  OAI211XLTS U3735 ( .A0(n4320), .A1(n12493), .B0(n4322), .C0(n4323), .Y(n4310) );
  NAND4XLTS U1985 ( .A(n2107), .B(n2439), .C(n2708), .D(n2709), .Y(n2707) );
  OAI211XLTS U1498 ( .A0(n11584), .A1(n10275), .B0(n1860), .C0(n1861), .Y(
        n1857) );
  OAI22XLTS U7322 ( .A0(n9491), .A1(n10061), .B0(n12356), .B1(n9845), .Y(n7647) );
  OAI211XLTS U6443 ( .A0(n9292), .A1(n11264), .B0(n6076), .C0(n6091), .Y(n6780) );
  OAI211XLTS U5930 ( .A0(n10512), .A1(n12400), .B0(n6476), .C0(n5361), .Y(
        n6472) );
  NAND4BXLTS U7183 ( .AN(n7353), .B(n7354), .C(n7355), .D(n7356), .Y(n7352) );
  OAI211XLTS U3675 ( .A0(n4224), .A1(n10389), .B0(n4225), .C0(n4226), .Y(n4213) );
  OAI211XLTS U5603 ( .A0(n11288), .A1(n12042), .B0(n6104), .C0(n5375), .Y(
        n6103) );
  OAI211XLTS U5798 ( .A0(n9402), .A1(n6338), .B0(n6339), .C0(n6340), .Y(n6336)
         );
  OAI31XLTS U6048 ( .A0(sa30[1]), .A1(n9966), .A2(n6583), .B0(n5308), .Y(n6582) );
  OAI211XLTS U5229 ( .A0(n10428), .A1(n11204), .B0(n5331), .C0(n5332), .Y(
        n5320) );
  NAND4XLTS U7129 ( .A(n7203), .B(n7204), .C(n7205), .D(n7206), .Y(n7202) );
  OAI211XLTS U2042 ( .A0(n2761), .A1(n11556), .B0(n2762), .C0(n2468), .Y(n2760) );
  OAI22XLTS U5824 ( .A0(n5769), .A1(n10484), .B0(n5660), .B1(n10976), .Y(n6377) );
  OAI211XLTS U4560 ( .A0(n9102), .A1(n11339), .B0(n4166), .C0(n4181), .Y(n4981) );
  OAI211XLTS U3972 ( .A0(n10425), .A1(n12444), .B0(n4604), .C0(n3524), .Y(
        n4600) );
  OAI211XLTS U7193 ( .A0(n10612), .A1(n11540), .B0(n7379), .C0(n7380), .Y(
        n7376) );
  NAND4BXLTS U5429 ( .AN(n5816), .B(n5817), .C(n5818), .D(n5819), .Y(n5772) );
  NAND4XLTS U3640 ( .A(n4171), .B(n4172), .C(n4173), .D(n4174), .Y(n4170) );
  OAI211XLTS U3916 ( .A0(n4304), .A1(n11713), .B0(n3631), .C0(n4535), .Y(n4534) );
  AOI32XLTS U3779 ( .A0(n10758), .A1(n4378), .A2(n9665), .B0(n9907), .B1(n4378), .Y(n4377) );
  NAND2XLTS U1809 ( .A(n2489), .B(n2490), .Y(n2488) );
  AOI32XLTS U5662 ( .A0(n10983), .A1(n6182), .A2(n9763), .B0(n10153), .B1(
        n6182), .Y(n6181) );
  OAI211XLTS U1901 ( .A0(n2617), .A1(n10288), .B0(n2618), .C0(n2227), .Y(n2616) );
  OAI211XLTS U7236 ( .A0(n7454), .A1(n9834), .B0(n7456), .C0(n7457), .Y(n7453)
         );
  NAND4XLTS U3731 ( .A(n4312), .B(n4313), .C(n4314), .D(n4315), .Y(n4311) );
  OAI211XLTS U7924 ( .A0(n7317), .A1(n10073), .B0(n8324), .C0(n8325), .Y(n8323) );
  NAND4XLTS U3668 ( .A(n4215), .B(n4216), .C(n4217), .D(n4218), .Y(n4214) );
  OAI211XLTS U1882 ( .A0(n2587), .A1(n10304), .B0(n2588), .C0(n2589), .Y(n2571) );
  NAND4XLTS U1867 ( .A(n1655), .B(n2573), .C(n2574), .D(n2575), .Y(n2572) );
  AOI211XLTS U5641 ( .A0(n5782), .A1(n6151), .B0(n5276), .C0(n6152), .Y(n6146)
         );
  OAI211XLTS U1654 ( .A0(n2216), .A1(n9720), .B0(n2218), .C0(n2219), .Y(n2215)
         );
  NAND4XLTS U5616 ( .A(n6125), .B(n6126), .C(n6127), .D(n6128), .Y(n6124) );
  OAI211XLTS U8669 ( .A0(n10041), .A1(n11539), .B0(n7803), .C0(n8647), .Y(
        n8629) );
  NAND4XLTS U2259 ( .A(n2203), .B(n1791), .C(n2972), .D(n2973), .Y(n2971) );
  NAND4XLTS U5588 ( .A(n6081), .B(n6082), .C(n6083), .D(n6084), .Y(n6080) );
  NAND4XLTS U8653 ( .A(n8642), .B(n8122), .C(n8643), .D(n7428), .Y(n8630) );
  OAI211XLTS U8066 ( .A0(n8441), .A1(n11109), .B0(n8442), .C0(n8280), .Y(n8440) );
  NAND4XLTS U4279 ( .A(n4359), .B(n3839), .C(n4880), .D(n4881), .Y(n4879) );
  OAI211XLTS U1813 ( .A0(n2499), .A1(n12097), .B0(n2500), .C0(n2501), .Y(n2498) );
  NAND4XLTS U1702 ( .A(n1831), .B(n1705), .C(n2301), .D(n2302), .Y(n2300) );
  OAI211XLTS U1828 ( .A0(n10008), .A1(n12555), .B0(n1792), .C0(n2522), .Y(
        n2521) );
  OAI211XLTS U3940 ( .A0(n4573), .A1(n11757), .B0(n4574), .C0(n4322), .Y(n4555) );
  NAND4XLTS U3930 ( .A(n4557), .B(n4558), .C(n4559), .D(n4560), .Y(n4556) );
  OAI31XLTS U3556 ( .A0(n9129), .A1(n4031), .A2(n9132), .B0(n3526), .Y(n4029)
         );
  OAI22XLTS U5671 ( .A0(n9287), .A1(n10189), .B0(n5639), .B1(n10417), .Y(n6188) );
  NAND4XLTS U1886 ( .A(n1654), .B(n2595), .C(n2596), .D(n2597), .Y(n2594) );
  OAI211XLTS U3527 ( .A0(n3977), .A1(n12549), .B0(n3978), .C0(n3979), .Y(n3976) );
  OAI31XLTS U3589 ( .A0(n9141), .A1(n4087), .A2(n9144), .B0(n3565), .Y(n4085)
         );
  NAND4XLTS U1667 ( .A(n1894), .B(n1743), .C(n2234), .D(n2235), .Y(n2233) );
  NAND4XLTS U3030 ( .A(n2044), .B(n2472), .C(n3292), .D(n3069), .Y(n3291) );
  NAND4XLTS U5635 ( .A(n6144), .B(n6145), .C(n6146), .D(n6147), .Y(n6143) );
  OAI31XLTS U5439 ( .A0(n9322), .A1(n5831), .A2(n9326), .B0(n5324), .Y(n5829)
         );
  NAND4XLTS U5508 ( .A(n5945), .B(n5946), .C(n5947), .D(n5948), .Y(n5944) );
  OAI211XLTS U3541 ( .A0(n9907), .A1(n12038), .B0(n4007), .C0(n4008), .Y(n4006) );
  NAND4BXLTS U7244 ( .AN(n7481), .B(n7482), .C(n7483), .D(n7484), .Y(n7480) );
  OAI211XLTS U8427 ( .A0(n9826), .A1(n12463), .B0(n8550), .C0(n7883), .Y(n8549) );
  OAI31XLTS U5472 ( .A0(n9339), .A1(n5887), .A2(n9533), .B0(n5363), .Y(n5885)
         );
  OAI211XLTS U5417 ( .A0(n10153), .A1(n11977), .B0(n5791), .C0(n5792), .Y(
        n5790) );
  NAND4XLTS U1601 ( .A(n2105), .B(n2106), .C(n2107), .D(n2108), .Y(n2104) );
  OAI22XLTS U5424 ( .A0(n9288), .A1(n10958), .B0(n9313), .B1(n12495), .Y(n5805) );
  AOI211XLTS U5813 ( .A0(n12063), .A1(n12281), .B0(n6365), .C0(n5571), .Y(
        n6363) );
  AOI211XLTS U7993 ( .A0(n12135), .A1(n8385), .B0(n8386), .C0(n8387), .Y(n8384) );
  OAI211XLTS U3785 ( .A0(n10938), .A1(n11708), .B0(n4380), .C0(n4381), .Y(
        n4366) );
  AOI31XLTS U7108 ( .A0(sa20[0]), .A1(n7154), .A2(n7155), .B0(n7156), .Y(n7153) );
  NAND4XLTS U3752 ( .A(n4341), .B(n4342), .C(n4343), .D(n4344), .Y(n4340) );
  OAI211XLTS U3333 ( .A0(n10164), .A1(n10943), .B0(n3488), .C0(n3489), .Y(
        n3485) );
  NAND4XLTS U4888 ( .A(n5079), .B(n5080), .C(n5081), .D(n5082), .Y(n5078) );
  OAI211XLTS U5213 ( .A0(n10413), .A1(n10818), .B0(n5286), .C0(n5287), .Y(
        n5283) );
  NAND4XLTS U7398 ( .A(n7203), .B(n7777), .C(n7778), .D(n7779), .Y(n7776) );
  NAND4XLTS U7992 ( .A(n8382), .B(n8383), .C(n8384), .D(n7574), .Y(n8381) );
  NAND4XLTS U5537 ( .A(n5817), .B(n5420), .C(n5999), .D(n6000), .Y(n5998) );
  NAND4BBXLTS U5812 ( .AN(n6361), .BN(n6362), .C(n6363), .D(n6364), .Y(n6360)
         );
  NAND4XLTS U3774 ( .A(n3489), .B(n4368), .C(n4369), .D(n4370), .Y(n4367) );
  NAND4BXLTS U3378 ( .AN(n3621), .B(n3622), .C(n3623), .D(n3624), .Y(n3602) );
  NAND3XLTS U3909 ( .A(n4526), .B(n4527), .C(n4528), .Y(n4525) );
  NAND4XLTS U7107 ( .A(n7151), .B(n7084), .C(n7152), .D(n7153), .Y(n7150) );
  OAI211XLTS U3721 ( .A0(n12414), .A1(n12380), .B0(n4290), .C0(n4291), .Y(
        n4289) );
  NAND4XLTS U5657 ( .A(n5287), .B(n6172), .C(n6173), .D(n6174), .Y(n6171) );
  AOI31XLTS U7139 ( .A0(n9860), .A1(n7226), .A2(n11076), .B0(n7228), .Y(n7225)
         );
  NAND4XLTS U3685 ( .A(n3970), .B(n3622), .C(n4232), .D(n4233), .Y(n4231) );
  NAND4XLTS U7835 ( .A(n8245), .B(n7954), .C(n8246), .D(n8247), .Y(n8244) );
  INVX1TS U6970 ( .A(n1284), .Y(n1287) );
  OAI211XLTS U1941 ( .A0(n9112), .A1(n10544), .B0(n2669), .C0(n2670), .Y(n1456) );
  INVX1TS U1321 ( .A(n1470), .Y(n1473) );
  NAND4XLTS U5227 ( .A(n5322), .B(n5323), .C(n5324), .D(n5325), .Y(n5321) );
  OAI211XLTS U5422 ( .A0(n5414), .A1(n12204), .B0(n5801), .C0(n5802), .Y(n5789) );
  NAND4XLTS U5238 ( .A(n5361), .B(n5362), .C(n5363), .D(n5364), .Y(n5360) );
  NAND4XLTS U3480 ( .A(n3877), .B(n3878), .C(n3879), .D(n3880), .Y(n3876) );
  NAND4XLTS U5374 ( .A(n5707), .B(n5708), .C(n5709), .D(n5710), .Y(n5706) );
  NAND4XLTS U3345 ( .A(n3524), .B(n3525), .C(n3526), .D(n3527), .Y(n3523) );
  NAND4XLTS U3356 ( .A(n3563), .B(n3564), .C(n3565), .D(n3566), .Y(n3562) );
  AOI2BB2XLTS U1338 ( .B0(n9489), .B1(n1565), .A0N(n1565), .A1N(n9490), .Y(
        N459) );
  AND4X1TS U3525 ( .A(n3604), .B(n3970), .C(n3971), .D(n3972), .Y(n1550) );
  CLKINVX2TS U8611 ( .A(n1565), .Y(n6997) );
  OAI211XLTS U1537 ( .A0(n9104), .A1(n12118), .B0(n1958), .C0(n1959), .Y(n1955) );
  CLKINVX2TS U7035 ( .A(n1560), .Y(n1558) );
  NAND4XLTS U2032 ( .A(n2742), .B(n2743), .C(n2132), .D(n2744), .Y(n2741) );
  NAND4XLTS U5362 ( .A(n5682), .B(n5683), .C(n5684), .D(n5685), .Y(n5681) );
  OAI211XLTS U5668 ( .A0(n10829), .A1(n11402), .B0(n6184), .C0(n6185), .Y(
        n6170) );
  INVX1TS U1700 ( .A(n1433), .Y(n1435) );
  INVX1TS U1330 ( .A(n1424), .Y(n1427) );
  NAND4XLTS U3373 ( .A(n3604), .B(n3605), .C(n3606), .D(n3607), .Y(n3603) );
  NAND4XLTS U7166 ( .A(n7305), .B(n7306), .C(n7307), .D(n7308), .Y(n7304) );
  CLKINVX2TS U1617 ( .A(n1344), .Y(n1341) );
  NAND2XLTS U7240 ( .A(n7468), .B(n7469), .Y(n7443) );
  AOI22XLTS U1353 ( .A0(n1588), .A1(n9309), .B0(n9310), .B1(n1590), .Y(N444)
         );
  NAND4XLTS U4860 ( .A(n4468), .B(n4286), .C(n3903), .D(n5061), .Y(n5060) );
  AOI22XLTS U1265 ( .A0(n1351), .A1(n9569), .B0(n9567), .B1(n1354), .Y(n1502)
         );
  AOI22XLTS U1345 ( .A0(n1574), .A1(n9394), .B0(n9395), .B1(n1576), .Y(N452)
         );
  NAND4XLTS U7544 ( .A(n7615), .B(n7957), .C(n7958), .D(n7959), .Y(n7956) );
  AOI22XLTS U1257 ( .A0(n1342), .A1(n9574), .B0(n9572), .B1(n1343), .Y(n1495)
         );
  OR4X2TS U5237 ( .A(n5357), .B(n5358), .C(n5359), .D(n5360), .Y(n5233) );
  INVX1TS U7500 ( .A(n6984), .Y(n1567) );
  OR4X2TS U3355 ( .A(n3559), .B(n3560), .C(n3561), .D(n3562), .Y(n3436) );
  NOR4XLTS U3479 ( .A(n3873), .B(n3874), .C(n3875), .D(n3876), .Y(n1594) );
  AOI22XLTS U1365 ( .A0(n1342), .A1(n9586), .B0(n9587), .B1(n1343), .Y(N435)
         );
  AOI22XLTS U1218 ( .A0(n1445), .A1(n9584), .B0(n9582), .B1(n1447), .Y(n1444)
         );
  INVX1TS U2225 ( .A(n1407), .Y(n1408) );
  AOI22XLTS U6969 ( .A0(n1284), .A1(n9514), .B0(n9512), .B1(n1287), .Y(n6958)
         );
  AOI22XLTS U1212 ( .A0(n1433), .A1(n9588), .B0(n9586), .B1(n1435), .Y(n1432)
         );
  AOI22XLTS U5128 ( .A0(n1574), .A1(n9410), .B0(n9408), .B1(n1576), .Y(n5211)
         );
  NAND4XLTS U7823 ( .A(n7468), .B(n8229), .C(n8230), .D(n7631), .Y(n8228) );
  NAND4BXLTS U3491 ( .AN(n3902), .B(n3903), .C(n3904), .D(n3905), .Y(n3901) );
  AOI22XLTS U7010 ( .A0(n6997), .A1(n9504), .B0(n9502), .B1(n1565), .Y(n6996)
         );
  AOI22XLTS U1327 ( .A0(n1433), .A1(n9572), .B0(n9573), .B1(n1435), .Y(N467)
         );
  AOI22XLTS U7033 ( .A0(n1558), .A1(n9495), .B0(n9493), .B1(n1560), .Y(n7017)
         );
  NAND4BXLTS U7318 ( .AN(n7633), .B(n7634), .C(n7306), .D(n7635), .Y(n1511) );
  AOI22XLTS U3247 ( .A0(n1588), .A1(n9325), .B0(n9323), .B1(n1590), .Y(n3414)
         );
  OR4X2TS U6353 ( .A(n6192), .B(n6078), .C(n6740), .D(n6741), .Y(n5175) );
  NAND4XLTS U3869 ( .A(n4468), .B(n4469), .C(n4470), .D(n4471), .Y(n4467) );
  OR4X2TS U4470 ( .A(n4389), .B(n4168), .C(n4941), .D(n4942), .Y(n3380) );
  OR4X2TS U7232 ( .A(n7442), .B(n7443), .C(n7444), .D(n7445), .Y(n1294) );
  AOI22XLTS U1164 ( .A0(n1341), .A1(n1342), .B0(n1343), .B1(n1344), .Y(n1334)
         );
  AOI22XLTS U1228 ( .A0(n1462), .A1(n9579), .B0(n9577), .B1(n1464), .Y(n1461)
         );
  NAND4XLTS U6743 ( .A(n6272), .B(n5977), .C(n5644), .D(n6859), .Y(n6858) );
  NAND4XLTS U5410 ( .A(n5402), .B(n5775), .C(n5776), .D(n5777), .Y(n5774) );
  INVX1TS U1332 ( .A(n1417), .Y(n1420) );
  CLKINVX2TS U1864 ( .A(n1397), .Y(n1396) );
  INVX1TS U3683 ( .A(n3372), .Y(n1549) );
  AOI22XLTS U1407 ( .A0(n1412), .A1(n9619), .B0(n9620), .B1(n1413), .Y(N400)
         );
  AOI22XLTS U7065 ( .A0(n1605), .A1(n1515), .B0(n1516), .B1(n1607), .Y(n7042)
         );
  AND4X1TS U5679 ( .A(n6081), .B(n5683), .C(n6060), .D(n6190), .Y(n1615) );
  AOI22XLTS U7018 ( .A0(n1563), .A1(n9499), .B0(n9497), .B1(n1562), .Y(n7006)
         );
  INVX1TS U1512 ( .A(n1486), .Y(n1310) );
  INVX1TS U5506 ( .A(n1771), .Y(n1773) );
  INVX1TS U4664 ( .A(n3433), .Y(n1583) );
  INVX1TS U7612 ( .A(n6933), .Y(n1608) );
  INVX1TS U5535 ( .A(n5166), .Y(n1534) );
  AOI2BB2XLTS U1341 ( .B0(w2[15]), .B1(n1568), .A0N(n1568), .A1N(w2[15]), .Y(
        N456) );
  INVX1TS U3906 ( .A(n1781), .Y(n1783) );
  AOI22XLTS U1293 ( .A0(n1470), .A1(n1407), .B0(n1408), .B1(n1473), .Y(n1526)
         );
  INVX1TS U6547 ( .A(n5230), .Y(n1569) );
  INVX1TS U5360 ( .A(n5247), .Y(n1622) );
  AOI22XLTS U1615 ( .A0(n1341), .A1(n9559), .B0(n9557), .B1(n1344), .Y(n2131)
         );
  AOI22XLTS U1190 ( .A0(n1399), .A1(n9592), .B0(n9590), .B1(n1401), .Y(n1393)
         );
  AOI22XLTS U1189 ( .A0(n1395), .A1(n1396), .B0(n1397), .B1(n1398), .Y(n1394)
         );
  AOI22XLTS U3504 ( .A0(n1993), .A1(n9301), .B0(n9299), .B1(n1995), .Y(n3935)
         );
  INVX1TS U7348 ( .A(n6935), .Y(n1528) );
  AOI22XLTS U1463 ( .A0(n1771), .A1(n9421), .B0(n9422), .B1(n1773), .Y(N388)
         );
  CLKINVX2TS U3330 ( .A(n1555), .Y(n3340) );
  AOI22XLTS U5072 ( .A0(n9149), .A1(n1771), .B0(n1773), .B1(n1618), .Y(n5146)
         );
  AOI22XLTS U1469 ( .A0(n1781), .A1(n9331), .B0(n9332), .B1(n1783), .Y(N382)
         );
  CLKINVX2TS U1906 ( .A(n1371), .Y(n1368) );
  AOI22XLTS U1379 ( .A0(n1612), .A1(n9404), .B0(n9405), .B1(n1614), .Y(N422)
         );
  AOI2BB2XLTS U1352 ( .B0(w0[10]), .B1(n1587), .A0N(n1587), .A1N(w0[10]), .Y(
        N445) );
  AOI2BB2XLTS U1318 ( .B0(w0[6]), .B1(n1555), .A0N(n1555), .A1N(w0[6]), .Y(
        N473) );
  AOI22XLTS U1244 ( .A0(n1424), .A1(n1486), .B0(n1310), .B1(n1427), .Y(n1485)
         );
  CLKINVX2TS U3832 ( .A(n1587), .Y(n3420) );
  AOI22XLTS U3905 ( .A0(n1781), .A1(n9291), .B0(n9289), .B1(n1783), .Y(n4523)
         );
  AOI22XLTS U7179 ( .A0(n7019), .A1(n1598), .B0(n1600), .B1(n9181), .Y(n7345)
         );
  AOI22XLTS U3298 ( .A0(n3372), .A1(n9311), .B0(n9309), .B1(n1549), .Y(n3460)
         );
  AOI2BB2XLTS U1344 ( .B0(w1[10]), .B1(n1573), .A0N(n1573), .A1N(w1[10]), .Y(
        N453) );
  AOI22XLTS U1547 ( .A0(n1993), .A1(n9340), .B0(n9341), .B1(n1995), .Y(N379)
         );
  AOI22XLTS U6968 ( .A0(n6960), .A1(n1515), .B0(n1516), .B1(n1601), .Y(n6959)
         );
  CLKINVX2TS U3307 ( .A(n1629), .Y(n3364) );
  AOI22XLTS U5179 ( .A0(n5166), .A1(n9396), .B0(n9394), .B1(n1534), .Y(n5258)
         );
  XOR2X1TS U2072 ( .A(n1462), .B(n9238), .Y(n1402) );
  INVX1TS U5788 ( .A(n1648), .Y(n1650) );
  AOI22XLTS U2028 ( .A0(n1385), .A1(n9550), .B0(n9548), .B1(n1388), .Y(n2739)
         );
  CLKINVX2TS U5714 ( .A(n1573), .Y(n5217) );
  AOI22XLTS U5193 ( .A0(n5230), .A1(n1612), .B0(n1614), .B1(n1569), .Y(n5269)
         );
  AOI22XLTS U3217 ( .A0(n1546), .A1(n9333), .B0(n9331), .B1(n1548), .Y(n3377)
         );
  XOR2X1TS U1450 ( .A(n1412), .B(n1315), .Y(n1361) );
  AOI22XLTS U3195 ( .A0(n1551), .A1(n9342), .B0(n9340), .B1(n1553), .Y(n3351)
         );
  INVX1TS U7043 ( .A(n6999), .Y(n7000) );
  AOI22XLTS U1170 ( .A0(n1355), .A1(n9606), .B0(n9604), .B1(n1357), .Y(n1349)
         );
  AOI22XLTS U1176 ( .A0(n1368), .A1(n1369), .B0(n1370), .B1(n1371), .Y(n1367)
         );
  AOI22XLTS U5121 ( .A0(n1577), .A1(n9414), .B0(n9412), .B1(n1579), .Y(n5202)
         );
  AOI22XLTS U5177 ( .A0(n5217), .A1(n9149), .B0(n1618), .B1(n1573), .Y(n5259)
         );
  AOI22XLTS U6961 ( .A0(n1273), .A1(n9519), .B0(n9517), .B1(n1275), .Y(n6948)
         );
  AOI22XLTS U6960 ( .A0(n1517), .A1(n1602), .B0(n1604), .B1(n1519), .Y(n6949)
         );
  AOI22XLTS U1131 ( .A0(n1273), .A1(n9470), .B0(n9468), .B1(n1275), .Y(n1272)
         );
  AOI22XLTS U1184 ( .A0(n1385), .A1(n1386), .B0(n9239), .B1(n1388), .Y(n1378)
         );
  INVX1TS U6973 ( .A(n1278), .Y(n1277) );
  AOI22XLTS U5157 ( .A0(n5196), .A1(n5123), .B0(n9146), .B1(n1580), .Y(n5242)
         );
  AOI22XLTS U3287 ( .A0(n1633), .A1(n1588), .B0(n1590), .B1(n1635), .Y(n3455)
         );
  AOI22XLTS U1250 ( .A0(n1329), .A1(n1355), .B0(n1357), .B1(n9257), .Y(n1490)
         );
  AOI22XLTS U1316 ( .A0(n1551), .A1(n9299), .B0(n9300), .B1(n1553), .Y(N475)
         );
  INVX1TS U5408 ( .A(n5159), .Y(n1535) );
  AOI22XLTS U5787 ( .A0(n1648), .A1(n9379), .B0(n9377), .B1(n1650), .Y(n6325)
         );
  AOI22XLTS U3306 ( .A0(n3364), .A1(n1546), .B0(n1548), .B1(n1629), .Y(n3465)
         );
  AOI22XLTS U7819 ( .A0(n1641), .A1(n9475), .B0(n9473), .B1(n1643), .Y(n8225)
         );
  CLKINVX2TS U5390 ( .A(n1776), .Y(n1774) );
  AOI22XLTS U7060 ( .A0(n6933), .A1(n1519), .B0(n1517), .B1(n1608), .Y(n7036)
         );
  AOI22XLTS U1413 ( .A0(n1641), .A1(n9517), .B0(n9518), .B1(n1643), .Y(N395)
         );
  AOI22XLTS U3240 ( .A0(n1591), .A1(n9329), .B0(n9327), .B1(n1593), .Y(n3405)
         );
  AOI22XLTS U1418 ( .A0(n1648), .A1(n9417), .B0(n9418), .B1(n1650), .Y(N390)
         );
  AOI22XLTS U5168 ( .A0(n1619), .A1(n1574), .B0(n1576), .B1(n1621), .Y(n5253)
         );
  CLKINVX2TS U7230 ( .A(n1513), .Y(n1512) );
  AOI22XLTS U3296 ( .A0(n3420), .A1(n9137), .B0(n1632), .B1(n1587), .Y(n3461)
         );
  AOI22XLTS U1313 ( .A0(n1546), .A1(n9289), .B0(n9290), .B1(n1548), .Y(N478)
         );
  XOR2X1TS U3949 ( .A(n9167), .B(n9140), .Y(n3381) );
  XOR2X1TS U3342 ( .A(n9101), .B(n9130), .Y(n3356) );
  AOI22XLTS U1303 ( .A0(n1536), .A1(n9385), .B0(n9386), .B1(n1538), .Y(N483)
         );
  AOI22XLTS U5095 ( .A0(n5174), .A1(n9271), .B0(n1611), .B1(n1647), .Y(n5173)
         );
  AOI22XLTS U3215 ( .A0(n3379), .A1(n9084), .B0(n1625), .B1(n1780), .Y(n3378)
         );
  INVX1TS U3681 ( .A(n3422), .Y(n3421) );
  AOI22XLTS U6944 ( .A0(n6923), .A1(n6924), .B0(n9155), .B1(n1645), .Y(n6922)
         );
  AOI22XLTS U5152 ( .A0(n5238), .A1(n5190), .B0(n9171), .B1(n9198), .Y(n5237)
         );
  AOI22XLTS U6985 ( .A0(n1512), .A1(n9509), .B0(n9507), .B1(n1513), .Y(n6970)
         );
  AOI22XLTS U3270 ( .A0(n3441), .A1(n3394), .B0(n9164), .B1(n9184), .Y(n3440)
         );
  CLKINVX2TS U1795 ( .A(n1353), .Y(n1352) );
  CLKINVX2TS U1575 ( .A(n1331), .Y(n1328) );
  XOR2X1TS U4191 ( .A(n9185), .B(n9100), .Y(n4024) );
  AOI22XLTS U5169 ( .A0(n5159), .A1(n9401), .B0(n9399), .B1(n1535), .Y(n5252)
         );
  XOR2X1TS U6074 ( .A(n9199), .B(n9117), .Y(n5824) );
  AOI22XLTS U1300 ( .A0(n1531), .A1(n9377), .B0(n9378), .B1(n1533), .Y(N486)
         );
  XOR2X1TS U2316 ( .A(n1480), .B(n1412), .Y(n2230) );
  AOI22XLTS U5388 ( .A0(n1774), .A1(n9387), .B0(n9385), .B1(n1776), .Y(n5732)
         );
  AOI22XLTS U5097 ( .A0(n1531), .A1(n9419), .B0(n9417), .B1(n1533), .Y(n5172)
         );
  AOI22XLTS U1256 ( .A0(n1445), .A1(n1372), .B0(n9247), .B1(n1447), .Y(n1496)
         );
  AOI22XLTS U5073 ( .A0(n1536), .A1(n9428), .B0(n9426), .B1(n1538), .Y(n5145)
         );
  AOI22XLTS U5163 ( .A0(n5247), .A1(n1538), .B0(n1536), .B1(n1622), .Y(n5246)
         );
  INVX1TS U3301 ( .A(n3416), .Y(n3415) );
  XNOR2X1TS U3466 ( .A(n10023), .B(n9133), .Y(n3345) );
  AOI22XLTS U3312 ( .A0(n3433), .A1(n1626), .B0(n1628), .B1(n1583), .Y(n3471)
         );
  AOI22XLTS U5194 ( .A0(n5182), .A1(n9391), .B0(n9389), .B1(n9209), .Y(n5268)
         );
  INVX1TS U7101 ( .A(n7007), .Y(n7008) );
  AOI22XLTS U3281 ( .A0(n3338), .A1(n1551), .B0(n1553), .B1(n9133), .Y(n3449)
         );
  AOI22XLTS U3314 ( .A0(n3386), .A1(n9306), .B0(n9304), .B1(n9194), .Y(n3470)
         );
  AOI22XLTS U5081 ( .A0(n5159), .A1(n9423), .B0(n9421), .B1(n1535), .Y(n5155)
         );
  XOR2X1TS U7424 ( .A(n1644), .B(n6943), .Y(n6991) );
  AOI22XLTS U7103 ( .A0(n6965), .A1(n9484), .B0(n9483), .B1(n9219), .Y(n7146)
         );
  AOI22XLTS U5187 ( .A0(n1615), .A1(n1531), .B0(n1533), .B1(n9768), .Y(n5263)
         );
  AOI22XLTS U5080 ( .A0(n5157), .A1(n1615), .B0(n9769), .B1(n1770), .Y(n5156)
         );
  INVX1TS U5172 ( .A(n5203), .Y(n5206) );
  INVX1TS U5533 ( .A(n5219), .Y(n5218) );
  CLKBUFX2TS U3317 ( .A(n3332), .Y(n3331) );
  AOI22XLTS U1158 ( .A0(n1328), .A1(n1329), .B0(n9257), .B1(n1331), .Y(n1321)
         );
  INVX1TS U5182 ( .A(n5213), .Y(n5212) );
  CLKBUFX2TS U5223 ( .A(n5150), .Y(n5147) );
  AOI2BB2XLTS U3182 ( .B0(n3335), .B1(n3336), .A0N(n3335), .A1N(n3336), .Y(
        n3334) );
  CLKBUFX2TS U5197 ( .A(n5126), .Y(n5125) );
  AOI22XLTS U1169 ( .A0(n1351), .A1(n1352), .B0(n1353), .B1(n1354), .Y(n1350)
         );
  AOI22XLTS U6978 ( .A0(n6965), .A1(n1598), .B0(n1600), .B1(n9219), .Y(n6964)
         );
  CLKBUFX2TS U1296 ( .A(n1317), .Y(n1316) );
  CLKBUFX2TS U7049 ( .A(n6953), .Y(n6950) );
  INVX1TS U1267 ( .A(n1449), .Y(n1448) );
  AOI2BB2XLTS U7344 ( .B0(n7023), .B1(n7703), .A0N(n7023), .A1N(n7703), .Y(
        n7702) );
  AOI2BB2XLTS U3746 ( .B0(n3363), .B1(n4338), .A0N(n3363), .A1N(n4338), .Y(
        n4337) );
  AOI2BB2XLTS U1309 ( .B0(n1395), .B1(n1544), .A0N(n1395), .A1N(n1544), .Y(
        n1543) );
  AOI2BB2XLTS U7565 ( .B0(n6932), .B1(n7996), .A0N(n6932), .A1N(n7996), .Y(
        n7995) );
  XNOR2X1TS U5252 ( .A(n9206), .B(n9753), .Y(n5197) );
  AOI22XLTS U6950 ( .A0(n6934), .A1(n6935), .B0(n1528), .B1(n6936), .Y(n6930)
         );
  CLKBUFX2TS U7253 ( .A(n6926), .Y(n6927) );
  AOI2BB2XLTS U7005 ( .B0(n6990), .B1(n9459), .A0N(n9459), .A1N(n6990), .Y(
        n6989) );
  AOI2BB2XLTS U6948 ( .B0(n6930), .B1(n6931), .A0N(n6930), .A1N(n6931), .Y(
        n6929) );
  AOI2BB2XLTS U5629 ( .B0(n5157), .B1(n6141), .A0N(n5157), .A1N(n6141), .Y(
        n6140) );
  AOI2BB2XLTS U1243 ( .B0(n1484), .B1(n1485), .A0N(n1484), .A1N(n1485), .Y(
        n1483) );
  AOI22XLTS U8032 ( .A0(n6951), .A1(n1276), .B0(n1279), .B1(n6952), .Y(n8223)
         );
  AOI2BB2XLTS U4189 ( .B0(n3379), .B1(n4800), .A0N(n3379), .A1N(n4800), .Y(
        n4799) );
  AOI2BB2XLTS U6072 ( .B0(n5174), .B1(n6600), .A0N(n5174), .A1N(n6600), .Y(
        n6599) );
  AOI22XLTS U5057 ( .A0(n5124), .A1(n9260), .B0(n12673), .B1(n9142), .Y(n5120)
         );
  AOI22XLTS U3227 ( .A0(n3390), .A1(n9074), .B0(n12674), .B1(n9100), .Y(n3389)
         );
  AOI2BB2XLTS U2314 ( .B0(n1399), .B1(n3018), .A0N(n1399), .A1N(n3018), .Y(
        n3017) );
  AOI2BB2XLTS U3445 ( .B0(n3337), .B1(n3808), .A0N(n3337), .A1N(n3808), .Y(
        n3807) );
  AOI2BB2XLTS U7422 ( .B0(n6923), .B1(n7807), .A0N(n6923), .A1N(n7807), .Y(
        n7806) );
  AOI22XLTS U5107 ( .A0(n5186), .A1(n9259), .B0(n5126), .B1(n9116), .Y(n5185)
         );
  AOI2BB2XLTS U5055 ( .B0(n5120), .B1(n5121), .A0N(n5120), .A1N(n5121), .Y(
        n5119) );
  AOI2BB2XLTS U5116 ( .B0(n5196), .B1(n9275), .A0N(n9275), .A1N(n5196), .Y(
        n5195) );
  AOI2BB2XLTS U5106 ( .B0(n5131), .B1(n5185), .A0N(n5131), .A1N(n5185), .Y(
        n5184) );
  AOI2BB2XLTS U3226 ( .B0(n12670), .B1(n3389), .A0N(n12670), .A1N(n3389), .Y(
        n3388) );
  AOI2BB2XLTS U3177 ( .B0(n3328), .B1(n3329), .A0N(n3328), .A1N(n3329), .Y(
        n3327) );
  OAI22XLTS U5124 ( .A0(n5207), .A1(n12763), .B0(n12686), .B1(n5208), .Y(N195)
         );
  AOI2BB2XLTS U5250 ( .B0(n5122), .B1(n5398), .A0N(n5122), .A1N(n5398), .Y(
        n5397) );
  AOI22XLTS U6945 ( .A0(n6925), .A1(n6926), .B0(n9794), .B1(n9151), .Y(n6921)
         );
  AOI2BB2XLTS U6943 ( .B0(n6921), .B1(n6922), .A0N(n6921), .A1N(n6922), .Y(
        n6920) );
  INVX1TS U5052 ( .A(sa00[5]), .Y(n5116) );
  AND2X2TS U4448 ( .A(n9892), .B(n10368), .Y(n4000) );
  AND2X2TS U5010 ( .A(n10318), .B(sa00[5]), .Y(n4806) );
  AND2X2TS U4457 ( .A(n9884), .B(n10743), .Y(n4785) );
  AND2X2TS U2565 ( .A(n9852), .B(sa32[1]), .Y(n2560) );
  AND2X2TS U5018 ( .A(n9278), .B(n9788), .Y(n4546) );
  AND2X2TS U6329 ( .A(n9816), .B(n10327), .Y(n5821) );
  AND2X2TS U6340 ( .A(n9808), .B(n10709), .Y(n6585) );
  AND2X2TS U2944 ( .A(sa10[2]), .B(n10700), .Y(n2429) );
  AND2X2TS U2746 ( .A(sa21[6]), .B(n9362), .Y(n2384) );
  AND2X2TS U2943 ( .A(sa10[6]), .B(n9282), .Y(n2428) );
  AND2X2TS U2747 ( .A(sa21[2]), .B(n10727), .Y(n2385) );
  OR3X1TS U6322 ( .A(n10716), .B(n9820), .C(n6728), .Y(n6040) );
  CLKINVX2TS U2917 ( .A(n3241), .Y(n3237) );
  CLKINVX2TS U2720 ( .A(n3181), .Y(n3177) );
  AND2X2TS U8390 ( .A(n8180), .B(n8540), .Y(n7967) );
  AND2X2TS U2532 ( .A(sa32[1]), .B(n3002), .Y(n2962) );
  CLKINVX2TS U8226 ( .A(n8468), .Y(n8022) );
  INVX2TS U1123 ( .A(n1262), .Y(n1258) );
  INVX1TS U8345 ( .A(n8523), .Y(n8414) );
  NAND2BX1TS U8569 ( .AN(n9571), .B(n8600), .Y(n7134) );
  OR3X1TS U5007 ( .A(n11163), .B(n10309), .C(n9237), .Y(n4807) );
  CLKINVX2TS U2767 ( .A(n3199), .Y(n2924) );
  CLKINVX2TS U2529 ( .A(n3001), .Y(n2998) );
  AND2X2TS U2519 ( .A(n3130), .B(n9063), .Y(n2563) );
  AND2X2TS U6915 ( .A(n6911), .B(n6319), .Y(n5733) );
  AND3X2TS U6874 ( .A(n9452), .B(sa01[4]), .C(n6674), .Y(n5574) );
  NAND2BX1TS U8755 ( .AN(n9581), .B(n8667), .Y(n7080) );
  CLKINVX2TS U6330 ( .A(n5625), .Y(n6534) );
  AND2X2TS U6936 ( .A(n6901), .B(n9392), .Y(n5959) );
  CLKINVX2TS U6337 ( .A(n6720), .Y(n6177) );
  CLKINVX2TS U2964 ( .A(n3259), .Y(n2848) );
  OR3X1TS U2570 ( .A(n3139), .B(n2036), .C(n10349), .Y(n2034) );
  OR3X1TS U2961 ( .A(sa10[0]), .B(sa10[3]), .C(n9716), .Y(n1945) );
  AND2X2TS U2550 ( .A(n2996), .B(n9048), .Y(n1663) );
  AND2X2TS U8710 ( .A(n9613), .B(n8648), .Y(n7208) );
  OR3X1TS U2764 ( .A(sa21[0]), .B(sa21[3]), .C(n9712), .Y(n1882) );
  AND2X2TS U4985 ( .A(n3925), .B(n5112), .Y(n3650) );
  AND2X2TS U4944 ( .A(n5103), .B(n9256), .Y(n3949) );
  AND2X2TS U4954 ( .A(n4334), .B(n5106), .Y(n3651) );
  NAND2X1TS U4082 ( .A(n11721), .B(n11225), .Y(n4712) );
  NOR2X1TS U7262 ( .A(n12560), .B(n11802), .Y(n7515) );
  NAND2XLTS U6813 ( .A(n10974), .B(n10474), .Y(n6655) );
  AND2X2TS U3134 ( .A(n9066), .B(n9684), .Y(n2650) );
  CLKBUFX2TS U6203 ( .A(n11668), .Y(n5415) );
  INVX1TS U4514 ( .A(n4632), .Y(n4964) );
  INVX1TS U4709 ( .A(n4704), .Y(n5022) );
  NAND2X1TS U8381 ( .A(n12171), .B(n11652), .Y(n8197) );
  NOR2XLTS U2614 ( .A(n11104), .B(n2319), .Y(n2392) );
  NAND3X1TS U7684 ( .A(n12082), .B(n11801), .C(n7134), .Y(n7250) );
  NAND2XLTS U2151 ( .A(n11152), .B(n11895), .Y(n2873) );
  NAND2XLTS U2076 ( .A(n11130), .B(n11870), .Y(n2797) );
  INVX1TS U6592 ( .A(n6504), .Y(n6821) );
  CLKINVX1TS U6812 ( .A(n6655), .Y(n6892) );
  AOI31X1TS U2065 ( .A0(sa03[1]), .A1(n9685), .A2(n11440), .B0(n2789), .Y(
        n2787) );
  NOR2XLTS U4686 ( .A(n4130), .B(n12216), .Y(n4205) );
  NAND2XLTS U4789 ( .A(n10827), .B(n12213), .Y(n4675) );
  NOR2XLTS U6569 ( .A(n10935), .B(n12271), .Y(n6115) );
  NOR2XLTS U6374 ( .A(n10908), .B(n12263), .Y(n6071) );
  AOI22X1TS U6779 ( .A0(n12056), .A1(n11330), .B0(n12300), .B1(n11742), .Y(
        n6882) );
  NOR2XLTS U4491 ( .A(n10831), .B(n12221), .Y(n4161) );
  AOI21X1TS U5295 ( .A0(n6456), .A1(n10920), .B0(n12426), .Y(n5510) );
  OAI22X1TS U7264 ( .A0(n10033), .A1(n11487), .B0(n12101), .B1(n11874), .Y(
        n7518) );
  AOI22X1TS U7621 ( .A0(n11457), .A1(n10623), .B0(n11082), .B1(n11078), .Y(
        n8045) );
  OAI22XLTS U4210 ( .A0(n4474), .A1(n10406), .B0(n12491), .B1(n9902), .Y(n4808) );
  NOR2X1TS U4922 ( .A(n11762), .B(n12491), .Y(n5094) );
  OAI22XLTS U4295 ( .A0(n4247), .A1(n9930), .B0(n11708), .B1(n10164), .Y(n4882) );
  OAI211X1TS U4593 ( .A0(n10845), .A1(n9916), .B0(n4992), .C0(n4603), .Y(n4990) );
  NAND2XLTS U7309 ( .A(n12625), .B(n10692), .Y(n7613) );
  OAI22X1TS U1502 ( .A0(n1868), .A1(n11147), .B0(n1725), .B1(n11900), .Y(n1867) );
  NOR2XLTS U6752 ( .A(n11348), .B(n11329), .Y(n6632) );
  INVX2TS U4511 ( .A(n3864), .Y(n3542) );
  OAI22X1TS U7675 ( .A0(n12100), .A1(n12077), .B0(n11114), .B1(n12463), .Y(
        n8091) );
  OAI211XLTS U4478 ( .A0(n4632), .A1(n10490), .B0(n4609), .C0(n4602), .Y(n4952) );
  OAI211XLTS U6361 ( .A0(n6432), .A1(n10428), .B0(n6409), .C0(n6402), .Y(n6751) );
  NAND2XLTS U4209 ( .A(n11769), .B(n9686), .Y(n4815) );
  INVX2TS U6394 ( .A(n5694), .Y(n5340) );
  NOR2XLTS U3939 ( .A(n11762), .B(n9675), .Y(n4572) );
  OAI22XLTS U2180 ( .A0(n10675), .A1(n11482), .B0(n10544), .B1(n10279), .Y(
        n2904) );
  OAI211X1TS U6476 ( .A0(n10898), .A1(n9946), .B0(n6791), .C0(n6403), .Y(n6789) );
  AOI22X1TS U5483 ( .A0(n10878), .A1(n11318), .B0(n11006), .B1(n11012), .Y(
        n5906) );
  OAI22X1TS U1526 ( .A0(n1931), .A1(n11126), .B0(n1763), .B1(n11877), .Y(n1930) );
  OAI211XLTS U6556 ( .A0(n6504), .A1(n10445), .B0(n6481), .C0(n6474), .Y(n6809) );
  OAI22X1TS U2105 ( .A0(n10662), .A1(n11472), .B0(n10570), .B1(n10255), .Y(
        n2828) );
  INVX2TS U3053 ( .A(n12288), .Y(n1991) );
  OAI211X1TS U6671 ( .A0(n10925), .A1(n9950), .B0(n6849), .C0(n6475), .Y(n6847) );
  AOI31XLTS U7945 ( .A0(n9898), .A1(n9366), .A2(n11897), .B0(n8342), .Y(n8336)
         );
  INVX2TS U2458 ( .A(n1807), .Y(n2577) );
  INVX2TS U6589 ( .A(n5719), .Y(n5379) );
  OAI22XLTS U2595 ( .A0(n2920), .A1(n12176), .B0(n1888), .B1(n1871), .Y(n3149)
         );
  OAI22X1TS U8283 ( .A0(n10346), .A1(n11647), .B0(n10097), .B1(n10357), .Y(
        n8515) );
  AOI22XLTS U3390 ( .A0(n11768), .A1(n10459), .B0(n10148), .B1(n11375), .Y(
        n3660) );
  INVX2TS U4706 ( .A(n3889), .Y(n3581) );
  NAND4X1TS U1989 ( .A(n2711), .B(n2712), .C(n2273), .D(n1903), .Y(n2710) );
  OAI211XLTS U4673 ( .A0(n4704), .A1(n10472), .B0(n4681), .C0(n4674), .Y(n5010) );
  AOI22X1TS U8050 ( .A0(n11916), .A1(n11928), .B0(n12369), .B1(n11156), .Y(
        n8432) );
  AOI22X1TS U5377 ( .A0(n10868), .A1(n5717), .B0(n10937), .B1(n12247), .Y(
        n5715) );
  OAI22X1TS U5772 ( .A0(n10173), .A1(n11753), .B0(n11372), .B1(n10225), .Y(
        n6305) );
  OAI22X1TS U1704 ( .A0(n2306), .A1(n12476), .B0(n10547), .B1(n10981), .Y(
        n2305) );
  OAI22X1TS U5491 ( .A0(n11366), .A1(n10919), .B0(n10511), .B1(n10217), .Y(
        n5911) );
  OAI22XLTS U5949 ( .A0(n5921), .A1(n10572), .B0(n9718), .B1(n10222), .Y(n6495) );
  AOI22XLTS U1839 ( .A0(n11506), .A1(n2217), .B0(n11953), .B1(n11052), .Y(
        n2538) );
  AOI221XLTS U5910 ( .A0(n5372), .A1(n9384), .B0(n11700), .B1(n11970), .C0(
        n6455), .Y(n6454) );
  OAI22X1TS U3755 ( .A0(n10788), .A1(n10939), .B0(n11804), .B1(n9908), .Y(
        n4346) );
  OAI211X1TS U2298 ( .A0(n11642), .A1(n12564), .B0(n3008), .C0(n3009), .Y(
        n3007) );
  OAI22X1TS U4307 ( .A0(n3615), .A1(n10754), .B0(n3616), .B1(n10789), .Y(n4891) );
  OAI22XLTS U2801 ( .A0(n2819), .A1(n11608), .B0(n12169), .B1(n11471), .Y(
        n3211) );
  OAI22XLTS U2952 ( .A0(n2297), .A1(n12468), .B0(n11465), .B1(n11600), .Y(
        n3253) );
  OAI211XLTS U7238 ( .A0(n11890), .A1(n11119), .B0(n7463), .C0(n7464), .Y(
        n7452) );
  OAI22XLTS U7982 ( .A0(n7466), .A1(n10750), .B0(n11176), .B1(n12128), .Y(
        n8375) );
  AOI31XLTS U6144 ( .A0(n11730), .A1(n10174), .A2(n10487), .B0(n9981), .Y(
        n6665) );
  OAI22X1TS U7794 ( .A0(n8190), .A1(n11166), .B0(n7465), .B1(n11641), .Y(n8185) );
  AOI22X1TS U3041 ( .A0(n10516), .A1(n12311), .B0(n12614), .B1(n12105), .Y(
        n3294) );
  AOI32X1TS U2237 ( .A0(n10000), .A1(n2956), .A2(n11947), .B0(n9721), .B1(
        n2956), .Y(n2955) );
  CLKINVX1TS U8027 ( .A(n8240), .Y(n8178) );
  OAI21X1TS U1937 ( .A0(n2059), .A1(n11853), .B0(n2667), .Y(n2666) );
  OAI31X1TS U2285 ( .A0(n12359), .A1(n12092), .A2(n12332), .B0(n11501), .Y(
        n2988) );
  OAI211X1TS U8163 ( .A0(n11108), .A1(n11597), .B0(n7823), .C0(n8284), .Y(
        n8474) );
  OAI22X1TS U7216 ( .A0(n7425), .A1(n9810), .B0(n7191), .B1(n11777), .Y(n7424)
         );
  OAI22X1TS U2119 ( .A0(n2246), .A1(n11465), .B0(n2815), .B1(n10219), .Y(n2840) );
  OAI211X1TS U1606 ( .A0(n2116), .A1(n11863), .B0(n2117), .C0(n2118), .Y(n2103) );
  NOR2XLTS U7365 ( .A(n11903), .B(n11109), .Y(n7717) );
  OAI211X1TS U2406 ( .A0(n12564), .A1(n9967), .B0(n3095), .C0(n1817), .Y(n3094) );
  OAI22X1TS U4180 ( .A0(n10789), .A1(n10502), .B0(n10944), .B1(n10922), .Y(
        n4797) );
  OAI22X1TS U4875 ( .A0(n12411), .A1(n10454), .B0(n11380), .B1(n10866), .Y(
        n5067) );
  INVX1TS U4933 ( .A(n3953), .Y(n4307) );
  OAI211XLTS U6169 ( .A0(n11690), .A1(n12205), .B0(n6686), .C0(n5822), .Y(
        n6683) );
  AOI22XLTS U1868 ( .A0(n12153), .A1(n11158), .B0(n12193), .B1(n10615), .Y(
        n2575) );
  OAI211X1TS U5694 ( .A0(n12385), .A1(n10892), .B0(n6208), .C0(n5453), .Y(
        n6205) );
  OAI22X1TS U2034 ( .A0(n10962), .A1(n11556), .B0(n10630), .B1(n12318), .Y(
        n2747) );
  OAI211X1TS U6215 ( .A0(n12211), .A1(n12496), .B0(n6709), .C0(n5802), .Y(
        n6708) );
  NAND2X1TS U2996 ( .A(n10235), .B(n11081), .Y(n2665) );
  INVX1TS U6005 ( .A(n5617), .Y(n5641) );
  CLKINVX2TS U5825 ( .A(n5995), .Y(n5660) );
  AOI22X1TS U6822 ( .A0(n10181), .A1(n5974), .B0(n10478), .B1(n6335), .Y(n6877) );
  OAI22X1TS U3494 ( .A0(n3913), .A1(n12533), .B0(n3914), .B1(n12381), .Y(n3908) );
  OAI22XLTS U7135 ( .A0(n7218), .A1(n12069), .B0(n11425), .B1(n10009), .Y(
        n7211) );
  AOI211X1TS U2280 ( .A0(n11520), .A1(n11058), .B0(n2992), .C0(n2993), .Y(
        n2990) );
  OAI211X1TS U6754 ( .A0(n11373), .A1(n10484), .B0(n6868), .C0(n6616), .Y(
        n6867) );
  OAI211XLTS U4871 ( .A0(n12206), .A1(n10871), .B0(n5070), .C0(n4818), .Y(
        n5069) );
  AOI22X1TS U3037 ( .A0(n11829), .A1(n3058), .B0(n11023), .B1(n2657), .Y(n3295) );
  OAI211X1TS U6497 ( .A0(n6195), .A1(n11359), .B0(n6795), .C0(n6796), .Y(n6794) );
  OAI22X1TS U8026 ( .A0(n8413), .A1(n10696), .B0(n8178), .B1(n12155), .Y(n8411) );
  INVX1TS U4122 ( .A(n3822), .Y(n3846) );
  AOI32X1TS U2322 ( .A0(n11062), .A1(n3025), .A2(n10192), .B0(n9923), .B1(
        n3025), .Y(n3024) );
  OAI22X1TS U4157 ( .A0(n9121), .A1(n10402), .B0(n12546), .B1(n11386), .Y(
        n4750) );
  OAI211X1TS U3860 ( .A0(n4459), .A1(n11256), .B0(n4460), .C0(n4461), .Y(n4458) );
  OAI211X1TS U1539 ( .A0(n1964), .A1(n11080), .B0(n1966), .C0(n1967), .Y(n1963) );
  AOI2BB2XLTS U3935 ( .B0(n12030), .B1(n4568), .A0N(n10775), .A1N(n9937), .Y(
        n4564) );
  OAI21X1TS U1719 ( .A0(n2339), .A1(n11905), .B0(n2340), .Y(n2337) );
  OAI211XLTS U8154 ( .A0(n9857), .A1(n11599), .B0(n8476), .C0(n7813), .Y(n8475) );
  OAI21X1TS U1684 ( .A0(n2272), .A1(n11881), .B0(n2273), .Y(n2270) );
  OAI211X1TS U2638 ( .A0(n11143), .A1(n1882), .B0(n3172), .C0(n1833), .Y(n3171) );
  OAI211X1TS U2410 ( .A0(n12562), .A1(n10292), .B0(n3008), .C0(n2545), .Y(
        n3093) );
  OAI211XLTS U5321 ( .A0(n5589), .A1(n11992), .B0(n5591), .C0(n5592), .Y(n5588) );
  AOI32X1TS U4739 ( .A0(n4432), .A1(n4207), .A2(n10388), .B0(n10810), .B1(
        n4207), .Y(n5026) );
  AOI32X1TS U4544 ( .A0(n4392), .A1(n4163), .A2(n10399), .B0(n10838), .B1(
        n4163), .Y(n4968) );
  AOI32X1TS U6427 ( .A0(n6195), .A1(n6073), .A2(n10526), .B0(n10903), .B1(
        n6073), .Y(n6767) );
  OAI21X1TS U1833 ( .A0(n2531), .A1(n11947), .B0(n2532), .Y(n2525) );
  OAI211XLTS U5474 ( .A0(n10920), .A1(n11307), .B0(n5893), .C0(n5894), .Y(
        n5892) );
  OAI211XLTS U3591 ( .A0(n10823), .A1(n11298), .B0(n4093), .C0(n4094), .Y(
        n4092) );
  OAI211X1TS U6663 ( .A0(n5928), .A1(n11216), .B0(n6846), .C0(n6507), .Y(n6845) );
  OAI211X1TS U4780 ( .A0(n4128), .A1(n11400), .B0(n5047), .C0(n4707), .Y(n5046) );
  OAI211X1TS U2419 ( .A0(n2552), .A1(n10175), .B0(n3096), .C0(n3097), .Y(n3085) );
  OAI211X1TS U6468 ( .A0(n5872), .A1(n11205), .B0(n6788), .C0(n6435), .Y(n6787) );
  OAI211XLTS U5240 ( .A0(n10445), .A1(n11216), .B0(n5370), .C0(n5371), .Y(
        n5359) );
  AOI211XLTS U3758 ( .A0(n3991), .A1(n4348), .B0(n3478), .C0(n4349), .Y(n4343)
         );
  OAI211X1TS U4585 ( .A0(n4072), .A1(n11411), .B0(n4989), .C0(n4635), .Y(n4988) );
  OAI211XLTS U3358 ( .A0(n10472), .A1(n11399), .B0(n3572), .C0(n3573), .Y(
        n3561) );
  AOI31X1TS U8065 ( .A0(n10340), .A1(n12370), .A2(n10078), .B0(n8440), .Y(
        n8439) );
  AOI211X1TS U7836 ( .A0(n12595), .A1(n7582), .B0(n7632), .C0(n8248), .Y(n8247) );
  NAND4X1TS U3482 ( .A(n3883), .B(n3884), .C(n3885), .D(n3886), .Y(n3882) );
  NAND4BX1TS U4132 ( .AN(n4009), .B(n3605), .C(n4752), .D(n4753), .Y(n4751) );
  NAND4X1TS U5364 ( .A(n5688), .B(n5689), .C(n5690), .D(n5691), .Y(n5687) );
  AND4X1TS U5290 ( .A(n5362), .B(n5495), .C(n5496), .D(n5497), .Y(n1581) );
  AND4X1TS U5265 ( .A(n5323), .B(n5429), .C(n5430), .D(n5431), .Y(n1623) );
  AND4X1TS U7191 ( .A(n7371), .B(n7151), .C(n7058), .D(n7372), .Y(n1557) );
  CLKINVX2TS U7180 ( .A(n1600), .Y(n1598) );
  INVX1TS U5599 ( .A(n1574), .Y(n1576) );
  INVX1TS U3651 ( .A(n1588), .Y(n1590) );
  CLKINVX2TS U8424 ( .A(n1607), .Y(n1605) );
  AND4X1TS U1452 ( .A(n1732), .B(n1733), .C(n1734), .D(n1735), .Y(n1318) );
  NAND4X1TS U1514 ( .A(n1732), .B(n1893), .C(n1894), .D(n1895), .Y(n1892) );
  AND4X1TS U2073 ( .A(n1893), .B(n1734), .C(n2792), .D(n2793), .Y(n1387) );
  AND4X1TS U1439 ( .A(n1694), .B(n1695), .C(n1696), .D(n1697), .Y(n1474) );
  AND4X1TS U7426 ( .A(n7677), .B(n7305), .C(n7808), .D(n7809), .Y(n1520) );
  AND4X1TS U2396 ( .A(n2595), .B(n2588), .C(n3083), .D(n3084), .Y(n1481) );
  INVX1TS U3505 ( .A(n1993), .Y(n1995) );
  AND4X1TS U1825 ( .A(n2204), .B(n2515), .C(n2516), .D(n2517), .Y(n1384) );
  AOI22XLTS U1337 ( .A0(n9485), .A1(n1562), .B0(n1563), .B1(n9483), .Y(N460)
         );
  AND4X1TS U3382 ( .A(n3631), .B(n3632), .C(n3633), .D(n3634), .Y(n1997) );
  INVX1TS U7136 ( .A(n6960), .Y(n1601) );
  INVX1TS U3750 ( .A(n1546), .Y(n1548) );
  AOI22XLTS U5056 ( .A0(n5122), .A1(n5123), .B0(n9145), .B1(n1778), .Y(n5121)
         );
  INVX1TS U5633 ( .A(n1531), .Y(n1533) );
  INVX1TS U1557 ( .A(n1355), .Y(n1357) );
  INVX1TS U3448 ( .A(n1551), .Y(n1553) );
  INVX1TS U5330 ( .A(n1536), .Y(n1538) );
  AND4X1TS U8036 ( .A(n8416), .B(n8417), .C(n8418), .D(n8419), .Y(n1529) );
  AOI22XLTS U3194 ( .A0(n9137), .A1(n1785), .B0(n1787), .B1(n1632), .Y(n3352)
         );
  AOI2BB2X1TS U1347 ( .B0(w1[13]), .B1(n1580), .A0N(n1580), .A1N(w1[13]), .Y(
        N450) );
  AOI22XLTS U1277 ( .A0(n1355), .A1(n9557), .B0(n9558), .B1(n1357), .Y(N499)
         );
  AOI22XLTS U1287 ( .A0(n1517), .A1(n9473), .B0(n9474), .B1(n1519), .Y(N491)
         );
  INVX1TS U5108 ( .A(n5133), .Y(n5131) );
  AOI22XLTS U1412 ( .A0(n1273), .A1(n9512), .B0(n9513), .B1(n1275), .Y(N396)
         );
  AOI22XLTS U1403 ( .A0(n1328), .A1(n9609), .B0(n9610), .B1(n1331), .Y(N402)
         );
  AOI22XLTS U7020 ( .A0(n1285), .A1(n7007), .B0(n7008), .B1(n1286), .Y(n7004)
         );
  AOI2BB2X1TS U7124 ( .B0(n1271), .B1(n7194), .A0N(n1271), .A1N(n7194), .Y(
        n7193) );
  INVX1TS U1251 ( .A(n1426), .Y(n1425) );
  AOI2BB2XLTS U5115 ( .B0(n5148), .B1(n5195), .A0N(n5148), .A1N(n5195), .Y(
        n5194) );
  AOI22X1TS U7036 ( .A0(n1303), .A1(n7018), .B0(n1282), .B1(n1304), .Y(n7015)
         );
  AOI2BB2XLTS U1198 ( .B0(n1323), .B1(n1411), .A0N(n1323), .A1N(n1411), .Y(
        n1410) );
  CLKINVX2TS U6938 ( .A(sa01[0]), .Y(n6917) );
  INVX2TS U6930 ( .A(sa01[4]), .Y(n6352) );
  NOR2X1TS U2780 ( .A(sa21[0]), .B(sa21[3]), .Y(n3191) );
  NOR2X1TS U8219 ( .A(sa31[0]), .B(sa31[3]), .Y(n8479) );
  NOR2X1TS U2977 ( .A(sa10[0]), .B(sa10[3]), .Y(n3251) );
  NOR3XLTS U5089 ( .A(n5167), .B(n11965), .C(dcnt[1]), .Y(N21) );
  CLKINVX2TS U4445 ( .A(n4742), .Y(n4922) );
  CLKAND2X2TS U8403 ( .A(n8271), .B(n8545), .Y(n7588) );
  CLKINVX2TS U6311 ( .A(n6738), .Y(n6048) );
  CLKAND2X2TS U8133 ( .A(n9898), .B(n9850), .Y(n7716) );
  NAND2XLTS U5890 ( .A(n11694), .B(n11408), .Y(n6440) );
  OAI22XLTS U7946 ( .A0(n7733), .A1(n10342), .B0(n10657), .B1(n10707), .Y(
        n8342) );
  NAND2X1TS U3997 ( .A(n10843), .B(n12406), .Y(n3862) );
  NAND3XLTS U7769 ( .A(n11426), .B(n11420), .C(n9802), .Y(n7178) );
  AOI22X1TS U2669 ( .A0(n12373), .A1(n11894), .B0(n11100), .B1(n11489), .Y(
        n3179) );
  AOI32XLTS U5239 ( .A0(sa23[0]), .A1(n10869), .A2(n5366), .B0(n10439), .B1(
        n10870), .Y(n5364) );
  AOI32XLTS U3357 ( .A0(n9840), .A1(n10901), .A2(n3568), .B0(n10475), .B1(
        n10900), .Y(n3566) );
  AOI22X1TS U2662 ( .A0(n11136), .A1(n1720), .B0(n12147), .B1(n9987), .Y(n3173) );
  AOI32XLTS U3346 ( .A0(sa11[0]), .A1(n10916), .A2(n3529), .B0(n10493), .B1(
        n10917), .Y(n3527) );
  AOI21XLTS U7416 ( .A0(n11832), .A1(n11437), .B0(n11766), .Y(n7791) );
  CLKINVX1TS U6397 ( .A(n6432), .Y(n6763) );
  OAI32X1TS U3994 ( .A0(sa11[6]), .A1(n9644), .A2(n11338), .B0(n4624), .B1(
        n10056), .Y(n3548) );
  AOI22X1TS U2433 ( .A0(n11058), .A1(n11596), .B0(n11453), .B1(n11913), .Y(
        n3106) );
  OAI222X1TS U7144 ( .A0(n11486), .A1(n11850), .B0(n12119), .B1(n12083), .C0(
        n10628), .C1(n9817), .Y(n7240) );
  AOI31X1TS U6156 ( .A0(n12681), .A1(n6674), .A2(n9974), .B0(n6675), .Y(n6667)
         );
  AOI21X1TS U5270 ( .A0(n10461), .A1(n10892), .B0(n12418), .Y(n5444) );
  OAI22XLTS U2792 ( .A0(n2844), .A1(n12169), .B0(n1951), .B1(n1934), .Y(n3209)
         );
  OAI22XLTS U2802 ( .A0(n11464), .A1(n12087), .B0(n11612), .B1(n10244), .Y(
        n3210) );
  OAI22XLTS U2605 ( .A0(n11476), .A1(n12079), .B0(n11631), .B1(n10268), .Y(
        n3150) );
  AOI22X1TS U5365 ( .A0(n10851), .A1(n5692), .B0(n5874), .B1(n12224), .Y(n5690) );
  OAI22X1TS U1524 ( .A0(n11602), .A1(n11608), .B0(n11121), .B1(n11614), .Y(
        n1919) );
  OAI22X1TS U1753 ( .A0(n2392), .A1(n10208), .B0(n10666), .B1(n12477), .Y(
        n2391) );
  OAI22X1TS U3608 ( .A0(n11254), .A1(n10822), .B0(n10419), .B1(n10114), .Y(
        n4111) );
  OAI21X1TS U7750 ( .A0(n11884), .A1(n11622), .B0(n11789), .Y(n8151) );
  AOI32X1TS U8431 ( .A0(n12321), .A1(n8556), .A2(n12083), .B0(n10681), .B1(
        n8556), .Y(n8553) );
  OAI211X1TS U6834 ( .A0(n11373), .A1(n10975), .B0(n6903), .C0(n6345), .Y(
        n6902) );
  AOI211X1TS U1493 ( .A0(n11941), .A1(n10284), .B0(n1842), .C0(n1843), .Y(
        n1839) );
  AOI22XLTS U7505 ( .A0(n11055), .A1(n11546), .B0(n12630), .B1(n12553), .Y(
        n7915) );
  OAI22XLTS U8505 ( .A0(n8057), .A1(n12464), .B0(n11487), .B1(n8061), .Y(n8589) );
  AOI22X1TS U2098 ( .A0(n12603), .A1(n9057), .B0(n11090), .B1(n10580), .Y(
        n2821) );
  OAI21X1TS U2408 ( .A0(n12192), .A1(n11913), .B0(n11918), .Y(n3095) );
  NOR2X1TS U6749 ( .A(n11355), .B(n10577), .Y(n5958) );
  OAI22X1TS U3459 ( .A0(n12284), .A1(n11386), .B0(n12039), .B1(n10124), .Y(
        n3832) );
  CLKINVX1TS U4356 ( .A(n4758), .Y(n4916) );
  OAI22X1TS U3783 ( .A0(n12547), .A1(n12038), .B0(n10108), .B1(n12064), .Y(
        n4375) );
  OAI22X1TS U5836 ( .A0(n9715), .A1(n12383), .B0(n9360), .B1(n11265), .Y(n6383) );
  OAI22XLTS U5828 ( .A0(n6378), .A1(n11373), .B0(n5668), .B1(n12021), .Y(n6358) );
  CLKINVX1TS U6238 ( .A(n6558), .Y(n6715) );
  NAND2XLTS U2251 ( .A(n9927), .B(n9964), .Y(n2224) );
  OAI22X1TS U5666 ( .A0(n12495), .A1(n11976), .B0(n10206), .B1(n12196), .Y(
        n6179) );
  AOI22XLTS U7095 ( .A0(n11037), .A1(n7128), .B0(n11444), .B1(n12088), .Y(
        n7115) );
  OAI21XLTS U7099 ( .A0(n12464), .A1(n12100), .B0(n7145), .Y(n7143) );
  OAI22X1TS U5428 ( .A0(n12204), .A1(n10206), .B0(n9965), .B1(n11689), .Y(
        n5815) );
  OAI22X1TS U2056 ( .A0(n2074), .A1(n11531), .B0(n11851), .B1(n11459), .Y(
        n2775) );
  AOI32X1TS U8520 ( .A0(n11486), .A1(n8063), .A2(n10678), .B0(n12337), .B1(
        n8063), .Y(n8597) );
  OAI22XLTS U5675 ( .A0(n6189), .A1(n10983), .B0(n5410), .B1(n10500), .Y(n6169) );
  AOI22X1TS U7130 ( .A0(n11065), .A1(n11782), .B0(n11433), .B1(n10590), .Y(
        n7204) );
  AOI22X1TS U3693 ( .A0(n10801), .A1(n4244), .B0(n10369), .B1(n4017), .Y(n4237) );
  OAI211X1TS U7417 ( .A0(n7798), .A1(n11604), .B0(n7800), .C0(n7801), .Y(n7790) );
  OAI31X1TS U7521 ( .A0(n11603), .A1(n9795), .A2(n9496), .B0(n7385), .Y(n7928)
         );
  OAI22XLTS U2755 ( .A0(n2364), .A1(n12484), .B0(n11477), .B1(n11618), .Y(
        n3193) );
  OAI22X1TS U5733 ( .A0(n11365), .A1(n10874), .B0(n10573), .B1(n10513), .Y(
        n6244) );
  OAI22XLTS U3793 ( .A0(n4386), .A1(n10757), .B0(n3612), .B1(n10787), .Y(n4365) );
  CLKINVX2TS U7921 ( .A(n8286), .Y(n7333) );
  OAI22XLTS U7185 ( .A0(n7119), .A1(n10033), .B0(n9825), .B1(n12084), .Y(n7351) );
  OAI22X1TS U5638 ( .A0(n10501), .A1(n10830), .B0(n11690), .B1(n10154), .Y(
        n6149) );
  AOI22X1TS U8287 ( .A0(n11497), .A1(n12134), .B0(n11171), .B1(n10691), .Y(
        n8519) );
  NAND4XLTS U4290 ( .A(n4769), .B(n4796), .C(n4268), .D(n4008), .Y(n4883) );
  OAI22XLTS U4880 ( .A0(n3962), .A1(n12381), .B0(n10872), .B1(n10867), .Y(
        n5072) );
  AOI211X1TS U4153 ( .A0(n10926), .A1(n11811), .B0(n4772), .C0(n4773), .Y(
        n4767) );
  OAI22X1TS U4553 ( .A0(n10109), .A1(n10398), .B0(n10486), .B1(n10850), .Y(
        n4978) );
  AOI211X1TS U8641 ( .A0(n11026), .A1(n10270), .B0(n8639), .C0(n7189), .Y(
        n8638) );
  OAI22XLTS U3946 ( .A0(n4578), .A1(n12206), .B0(n3910), .B1(n12573), .Y(n4554) );
  OAI211XLTS U4202 ( .A0(n12023), .A1(n11756), .B0(n4813), .C0(n4331), .Y(
        n4810) );
  AOI32XLTS U8074 ( .A0(n10724), .A1(n8450), .A2(n11529), .B0(n11557), .B1(
        n8450), .Y(n8449) );
  OAI211X1TS U4743 ( .A0(n4099), .A1(n10131), .B0(n4722), .C0(n3573), .Y(n5037) );
  AOI211X1TS U2838 ( .A0(n10557), .A1(n9057), .B0(n1918), .C0(n2827), .Y(n3232) );
  OAI21XLTS U8464 ( .A0(n7365), .A1(n10329), .B0(n8043), .Y(n8576) );
  NAND4XLTS U8626 ( .A(n7381), .B(n8625), .C(n8626), .D(n8627), .Y(n8615) );
  AOI22X1TS U2364 ( .A0(n11815), .A1(n2642), .B0(n10587), .B1(n2470), .Y(n3055) );
  OAI22XLTS U3873 ( .A0(n4319), .A1(n11381), .B0(n4297), .B1(n11756), .Y(n4472) );
  AOI211X1TS U2284 ( .A0(n11518), .A1(n10680), .B0(n2994), .C0(n2995), .Y(
        n2989) );
  OAI211X1TS U5719 ( .A0(n5899), .A1(n10918), .B0(n6239), .C0(n6240), .Y(n6238) );
  OAI22XLTS U4066 ( .A0(n4121), .A1(n10372), .B0(n9654), .B1(n10118), .Y(n4695) );
  AOI22X1TS U1956 ( .A0(n10552), .A1(n9065), .B0(n11893), .B1(n2686), .Y(n2684) );
  AOI211XLTS U3669 ( .A0(n12579), .A1(n9643), .B0(n4219), .C0(n4220), .Y(n4218) );
  AOI211X1TS U4384 ( .A0(n10369), .A1(n10430), .B0(n4930), .C0(n4263), .Y(
        n4927) );
  OAI211X1TS U7394 ( .A0(n7766), .A1(n11933), .B0(n7768), .C0(n7769), .Y(n7758) );
  AOI22X1TS U4337 ( .A0(n11799), .A1(n4780), .B0(n10122), .B1(n3992), .Y(n4910) );
  OAI211X1TS U4548 ( .A0(n4043), .A1(n10139), .B0(n4650), .C0(n3534), .Y(n4979) );
  OAI22X1TS U3991 ( .A0(n4065), .A1(n10377), .B0(n9658), .B1(n10110), .Y(n4623) );
  AOI31X1TS U4094 ( .A0(n4197), .A1(n10080), .A2(n10128), .B0(n4452), .Y(n4719) );
  CLKINVX2TS U2435 ( .A(n2222), .Y(n2038) );
  OAI211XLTS U8003 ( .A0(n11182), .A1(n10744), .B0(n8388), .C0(n8389), .Y(
        n8380) );
  OAI22X1TS U5874 ( .A0(n5865), .A1(n10567), .B0(n9714), .B1(n10214), .Y(n6423) );
  AOI22XLTS U2249 ( .A0(n10172), .A1(n2224), .B0(n12359), .B1(n2619), .Y(n2957) );
  AOI221X1TS U3952 ( .A0(n3535), .A1(n9183), .B0(n11751), .B1(n12057), .C0(
        n4583), .Y(n4582) );
  CLKINVX1TS U3944 ( .A(n3927), .Y(n4304) );
  AOI211X1TS U7619 ( .A0(n8047), .A1(n10735), .B0(n8048), .C0(n8049), .Y(n8046) );
  OAI22XLTS U7757 ( .A0(n7406), .A1(n11604), .B0(n7802), .B1(n7185), .Y(n8155)
         );
  OAI22XLTS U4267 ( .A0(n3953), .A1(n12530), .B0(n3917), .B1(n9651), .Y(n4868)
         );
  OAI211X1TS U6626 ( .A0(n5899), .A1(n10165), .B0(n6522), .C0(n5371), .Y(n6836) );
  AOI22XLTS U7199 ( .A0(n11878), .A1(n7074), .B0(n11885), .B1(n7394), .Y(n7387) );
  AOI22X1TS U1499 ( .A0(n12601), .A1(n11577), .B0(n10271), .B1(n1864), .Y(
        n1861) );
  OAI211X1TS U1492 ( .A0(n11906), .A1(n11901), .B0(n1839), .C0(n1840), .Y(
        n1836) );
  OAI211X1TS U6431 ( .A0(n5843), .A1(n10157), .B0(n6450), .C0(n5332), .Y(n6778) );
  OAI22XLTS U7279 ( .A0(n7549), .A1(n10328), .B0(n7246), .B1(n12334), .Y(n7540) );
  AOI211X1TS U6038 ( .A0(n10246), .A1(n11981), .B0(n6574), .C0(n6575), .Y(
        n6566) );
  AOI22XLTS U4241 ( .A0(n11213), .A1(n4850), .B0(n11249), .B1(n4324), .Y(n4848) );
  OAI211X1TS U2912 ( .A0(n12458), .A1(n11876), .B0(n3256), .C0(n3257), .Y(
        n3255) );
  OAI211XLTS U1954 ( .A0(n12175), .A1(n11626), .B0(n2684), .C0(n2685), .Y(
        n2683) );
  NAND4X1TS U6784 ( .A(n6610), .B(n6888), .C(n6889), .D(n6620), .Y(n6886) );
  AOI32X1TS U5692 ( .A0(n11253), .A1(n6207), .A2(n10436), .B0(n10566), .B1(
        n6207), .Y(n6206) );
  OAI211X1TS U5540 ( .A0(n9356), .A1(n10957), .B0(n6004), .C0(n6005), .Y(n6002) );
  AOI211X1TS U2044 ( .A0(n12338), .A1(n10519), .B0(n2763), .C0(n2764), .Y(
        n2762) );
  NAND4XLTS U7197 ( .A(n7386), .B(n7387), .C(n7388), .D(n7389), .Y(n7374) );
  OAI22XLTS U3548 ( .A0(n3628), .A1(n10794), .B0(n9122), .B1(n12548), .Y(n4019) );
  OAI22XLTS U3728 ( .A0(n9938), .A1(n12531), .B0(n4304), .B1(n10783), .Y(n4302) );
  OAI211X1TS U3688 ( .A0(n9169), .A1(n10793), .B0(n4237), .C0(n4238), .Y(n4235) );
  OAI22X1TS U3532 ( .A0(n3616), .A1(n10763), .B0(n3618), .B1(n10124), .Y(n3974) );
  OAI22XLTS U3739 ( .A0(n3914), .A1(n11715), .B0(n3916), .B1(n9651), .Y(n4308)
         );
  AOI32XLTS U5844 ( .A0(n6393), .A1(n11203), .A2(n11252), .B0(n10213), .B1(
        n6393), .Y(n6392) );
  OAI211X1TS U4333 ( .A0(n3841), .A1(n12548), .B0(n4910), .C0(n4016), .Y(n4909) );
  AOI31X1TS U8471 ( .A0(n9829), .A1(n12102), .A2(n12307), .B0(n7106), .Y(n8577) );
  OAI211X1TS U2430 ( .A0(n2038), .A1(n9999), .B0(n3106), .C0(n3107), .Y(n3105)
         );
  OAI211X1TS U2835 ( .A0(n11121), .A1(n1945), .B0(n3232), .C0(n1896), .Y(n3231) );
  AOI31X1TS U2383 ( .A0(n9526), .A1(n9059), .A2(n9688), .B0(n3076), .Y(n3073)
         );
  OAI211XLTS U7326 ( .A0(n7659), .A1(n11527), .B0(n7660), .C0(n7661), .Y(n7638) );
  AOI32X1TS U6622 ( .A0(n6235), .A1(n6117), .A2(n10535), .B0(n10930), .B1(
        n6117), .Y(n6825) );
  OAI211X1TS U6604 ( .A0(n10217), .A1(n10452), .B0(n6830), .C0(n6831), .Y(
        n6829) );
  AOI22X1TS U7655 ( .A0(n10733), .A1(n12313), .B0(n10257), .B1(n7121), .Y(
        n8078) );
  OAI211X1TS U2382 ( .A0(n3035), .A1(n11532), .B0(n3073), .C0(n3074), .Y(n3072) );
  OAI211XLTS U5822 ( .A0(n6374), .A1(n12004), .B0(n5961), .C0(n6375), .Y(n6359) );
  AOI211X1TS U2861 ( .A0(n11085), .A1(n11870), .B0(n2414), .C0(n2433), .Y(
        n3238) );
  OAI211X1TS U7654 ( .A0(n11113), .A1(n10329), .B0(n8077), .C0(n8078), .Y(
        n8076) );
  OAI211X1TS U3347 ( .A0(n10490), .A1(n11412), .B0(n3533), .C0(n3534), .Y(
        n3522) );
  OAI211XLTS U3880 ( .A0(n9902), .A1(n11382), .B0(n4484), .C0(n4485), .Y(n4328) );
  OAI211X1TS U4305 ( .A0(n3512), .A1(n9908), .B0(n4341), .C0(n4890), .Y(n4878)
         );
  AOI211X1TS U3931 ( .A0(n10390), .A1(n11212), .B0(n4561), .C0(n3654), .Y(
        n4558) );
  AOI211X1TS U2664 ( .A0(n11100), .A1(n11894), .B0(n2370), .C0(n2389), .Y(
        n3178) );
  AOI32X1TS U8548 ( .A0(n7890), .A1(n8604), .A2(n12558), .B0(n12077), .B1(
        n8604), .Y(n7861) );
  AOI211X1TS U7213 ( .A0(n10289), .A1(n12109), .B0(n7419), .C0(n7044), .Y(
        n7415) );
  NAND4XLTS U7614 ( .A(n8038), .B(n7562), .C(n8039), .D(n7506), .Y(n8037) );
  OAI211XLTS U3546 ( .A0(n3616), .A1(n12283), .B0(n4015), .C0(n4016), .Y(n4005) );
  OAI211X1TS U4522 ( .A0(n3722), .A1(n12405), .B0(n4970), .C0(n4646), .Y(n4969) );
  OAI211X1TS U6405 ( .A0(n5477), .A1(n12416), .B0(n6769), .C0(n6446), .Y(n6768) );
  NAND4XLTS U7698 ( .A(n8104), .B(n7379), .C(n8105), .D(n7413), .Y(n8103) );
  OAI211XLTS U8303 ( .A0(n8408), .A1(n11183), .B0(n8524), .C0(n7574), .Y(n8511) );
  OAI211X1TS U4717 ( .A0(n3788), .A1(n12395), .B0(n5028), .C0(n4718), .Y(n5027) );
  NAND4BXLTS U5260 ( .AN(n5419), .B(n5420), .C(n5421), .D(n5422), .Y(n5400) );
  NAND4X1TS U7209 ( .A(n7413), .B(n7414), .C(n7415), .D(n7083), .Y(n7412) );
  OAI211X1TS U6600 ( .A0(n5543), .A1(n12424), .B0(n6827), .C0(n6518), .Y(n6826) );
  NAND4BX1TS U6015 ( .AN(n5793), .B(n5403), .C(n6552), .D(n6553), .Y(n6551) );
  NAND4XLTS U5255 ( .A(n5402), .B(n5403), .C(n5404), .D(n5405), .Y(n5401) );
  AOI2BB2XLTS U1377 ( .B0(w2[23]), .B1(n9151), .A0N(n9152), .A1N(w2[23]), .Y(
        N424) );
  NOR4XLTS U6076 ( .A(n5562), .B(n6601), .C(n6602), .D(n6603), .Y(n5186) );
  AOI22XLTS U1325 ( .A0(n1445), .A1(n9567), .B0(n9568), .B1(n1447), .Y(N468)
         );
  AOI22XLTS U1363 ( .A0(n1351), .A1(n9582), .B0(n9583), .B1(n1354), .Y(N436)
         );
  AOI2BB2XLTS U1339 ( .B0(w2[13]), .B1(n1566), .A0N(n1566), .A1N(w2[13]), .Y(
        N458) );
  AOI22XLTS U1285 ( .A0(n1515), .A1(n9468), .B0(n9469), .B1(n1516), .Y(N492)
         );
  AOI22XLTS U1374 ( .A0(n1605), .A1(n9502), .B0(n9503), .B1(n1607), .Y(N427)
         );
  NAND4BX1TS U5211 ( .AN(n5276), .B(n5277), .C(n5278), .D(n5279), .Y(n1540) );
  AOI2BB2XLTS U1467 ( .B0(w1[31]), .B1(n9116), .A0N(n9117), .A1N(w1[31]), .Y(
        N384) );
  AOI22XLTS U1373 ( .A0(n1602), .A1(n9497), .B0(n9498), .B1(n1604), .Y(N428)
         );
  AOI22XLTS U1322 ( .A0(n1462), .A1(n9562), .B0(n9563), .B1(n1464), .Y(N470)
         );
  OAI211X1TS U1983 ( .A0(n9108), .A1(n2262), .B0(n2702), .C0(n2703), .Y(n1370)
         );
  AOI22XLTS U1401 ( .A0(n1341), .A1(n9604), .B0(n9605), .B1(n1344), .Y(N403)
         );
  AOI2BB2XLTS U1470 ( .B0(w0[26]), .B1(n1784), .A0N(n1784), .A1N(w0[26]), .Y(
        N381) );
  AOI22XLTS U1354 ( .A0(n1591), .A1(n9314), .B0(n9315), .B1(n1593), .Y(N443)
         );
  XNOR2XLTS U7126 ( .A(n1512), .B(n1560), .Y(n7195) );
  INVX1TS U7949 ( .A(n1273), .Y(n1275) );
  AOI22XLTS U1346 ( .A0(n1577), .A1(n9399), .B0(n9400), .B1(n1579), .Y(N451)
         );
  CLKINVX2TS U7001 ( .A(n6942), .Y(n6941) );
  AOI2BB2XLTS U1468 ( .B0(w0[24]), .B1(n1780), .A0N(n1780), .A1N(w0[24]), .Y(
        N383) );
  AOI2BB2XLTS U3184 ( .B0(n3339), .B1(n3340), .A0N(n3340), .A1N(n3339), .Y(
        n3335) );
  INVX1TS U6996 ( .A(n6936), .Y(n6934) );
  AOI22XLTS U1397 ( .A0(n1368), .A1(n9594), .B0(n9595), .B1(n1371), .Y(N405)
         );
  AOI2BB2XLTS U1416 ( .B0(w2[31]), .B1(n9127), .A0N(n9128), .A1N(w2[31]), .Y(
        N392) );
  AOI2BB2XLTS U1414 ( .B0(w2[29]), .B1(n1644), .A0N(n1644), .A1N(w2[29]), .Y(
        N394) );
  CLKINVX1TS U7021 ( .A(n1286), .Y(n1285) );
  CLKINVX1TS U3291 ( .A(n3409), .Y(n3406) );
  AOI22X1TS U3242 ( .A0(n3406), .A1(n3407), .B0(n3408), .B1(n3409), .Y(n3403)
         );
  AOI22XLTS U5142 ( .A0(n5225), .A1(n5204), .B0(n5205), .B1(n5226), .Y(n5222)
         );
  AOI22X1TS U1213 ( .A0(n1436), .A1(n1437), .B0(n1438), .B1(n1439), .Y(n1430)
         );
  AOI22X1TS U1276 ( .A0(n1369), .A1(n1397), .B0(n1396), .B1(n9251), .Y(n1509)
         );
  AOI22XLTS U7013 ( .A0(n6998), .A1(n6999), .B0(n7000), .B1(n7001), .Y(n6994)
         );
  AOI22XLTS U1199 ( .A0(n1412), .A1(n9269), .B0(n1317), .B1(n1413), .Y(n1411)
         );
  NOR4XLTS U8798 ( .A(n5318), .B(n5319), .C(n5320), .D(n5321), .Y(n5124) );
  NOR4XLTS U8799 ( .A(n7704), .B(n7705), .C(n7706), .D(n7707), .Y(n6935) );
  NOR4XLTS U8800 ( .A(n3482), .B(n4877), .C(n4878), .D(n4879), .Y(n3441) );
  NOR4XLTS U8801 ( .A(n3520), .B(n3521), .C(n3522), .D(n3523), .Y(n3330) );
  NOR4XLTS U8802 ( .A(n5771), .B(n5772), .C(n5773), .D(n5774), .Y(n5159) );
  NOR4XLTS U8803 ( .A(n2207), .B(n1813), .C(n2519), .D(n2944), .Y(n1407) );
  NOR4XLTS U8804 ( .A(n2101), .B(n2102), .C(n2103), .D(n2104), .Y(n1329) );
  AOI21X1TS U8805 ( .A0(n12206), .A1(n11773), .B0(n12490), .Y(n8680) );
  OA22X1TS U8806 ( .A0(n12490), .A1(n9639), .B0(n12538), .B1(n10406), .Y(n8681) );
  NAND4X1TS U8807 ( .A(n4874), .B(n4822), .C(n4814), .D(n8681), .Y(n8682) );
  AOI211X1TS U8808 ( .A0(n11374), .A1(n10814), .B0(n8680), .C0(n8682), .Y(
        n8683) );
  AOI211X1TS U8809 ( .A0(n12201), .A1(n10115), .B0(n4832), .C0(n4566), .Y(
        n8684) );
  OAI211X1TS U8810 ( .A0(n4319), .A1(n12379), .B0(n8683), .C0(n8684), .Y(n4292) );
  OAI211X1TS U8811 ( .A0(n9711), .A1(n12012), .B0(n6620), .C0(n6285), .Y(n8685) );
  AOI21X1TS U8812 ( .A0(n10237), .A1(n6617), .B0(n8685), .Y(n8686) );
  OAI211X1TS U8813 ( .A0(n10174), .A1(n10234), .B0(n6616), .C0(n8686), .Y(
        n8687) );
  AOI21X1TS U8814 ( .A0(n10549), .A1(n6306), .B0(n8687), .Y(n6353) );
  NAND4BX1TS U8815 ( .AN(n9749), .B(n12564), .C(n10287), .D(n1824), .Y(n8688)
         );
  AOI22X1TS U8816 ( .A0(n11911), .A1(n12151), .B0(n1820), .B1(n12358), .Y(
        n8689) );
  OAI211X1TS U8817 ( .A0(n10292), .A1(n9995), .B0(n8689), .C0(n1817), .Y(n8690) );
  AOI211X1TS U8818 ( .A0(n11918), .A1(n8688), .B0(n1813), .C0(n8690), .Y(n8691) );
  AOI22X1TS U8819 ( .A0(n11596), .A1(n1806), .B0(n1802), .B1(n12648), .Y(n8692) );
  OAI211X1TS U8820 ( .A0(n1689), .A1(n1804), .B0(n1799), .C0(n8692), .Y(n8693)
         );
  OAI22X1TS U8821 ( .A0(n1807), .A1(n9999), .B0(n1809), .B1(n11588), .Y(n8694)
         );
  NOR4XLTS U8822 ( .A(n1795), .B(n1796), .C(n8693), .D(n8694), .Y(n8695) );
  AND4X1TS U8823 ( .A(n1791), .B(n8691), .C(n1792), .D(n8695), .Y(n1340) );
  OAI22X1TS U8824 ( .A0(n7275), .A1(n11951), .B0(n10356), .B1(n11646), .Y(
        n8696) );
  AOI22X1TS U8825 ( .A0(n11192), .A1(n12597), .B0(n10310), .B1(n8219), .Y(
        n8697) );
  OAI21X1TS U8826 ( .A0(n9834), .A1(n10745), .B0(n8697), .Y(n8698) );
  AOI211X1TS U8827 ( .A0(n11170), .A1(n11503), .B0(n8696), .C0(n8698), .Y(
        n7616) );
  OAI22X1TS U8828 ( .A0(n5641), .A1(n9941), .B0(n5639), .B1(n10958), .Y(n8699)
         );
  AOI21X1TS U8829 ( .A0(n11208), .A1(n6187), .B0(n8699), .Y(n8700) );
  OAI22X1TS U8830 ( .A0(n6544), .A1(n12205), .B0(n6189), .B1(n12439), .Y(n8701) );
  AO22X1TS U8831 ( .A0(n10246), .A1(n5614), .B0(n5779), .B1(n12448), .Y(n8702)
         );
  AOI211X1TS U8832 ( .A0(n10840), .A1(n9969), .B0(n8701), .C0(n8702), .Y(n8703) );
  OAI211X1TS U8833 ( .A0(n9313), .A1(n10501), .B0(n8700), .C0(n8703), .Y(n8704) );
  AOI22X1TS U8834 ( .A0(n10563), .A1(n10142), .B0(n10496), .B1(n9283), .Y(
        n8705) );
  OAI211X1TS U8835 ( .A0(n11978), .A1(n10991), .B0(n5811), .C0(n5802), .Y(
        n8706) );
  OAI31X1TS U8836 ( .A0(sa30[2]), .A1(n6534), .A2(n12197), .B0(n6173), .Y(
        n8707) );
  OAI22X1TS U8837 ( .A0(n12496), .A1(n12440), .B0(n11403), .B1(n10150), .Y(
        n8708) );
  NOR4XLTS U8838 ( .A(n5814), .B(n8706), .C(n8707), .D(n8708), .Y(n8709) );
  NAND4BX1TS U8839 ( .AN(n8704), .B(n8705), .C(n5404), .D(n8709), .Y(n8710) );
  NOR3X1TS U8840 ( .A(n5787), .B(n5997), .C(n8710), .Y(n5182) );
  OAI211X1TS U8841 ( .A0(n10406), .A1(n12379), .B0(n4822), .C0(n4496), .Y(
        n8711) );
  AOI21X1TS U8842 ( .A0(n9189), .A1(n4819), .B0(n8711), .Y(n8712) );
  OAI211X1TS U8843 ( .A0(n10859), .A1(n11761), .B0(n4818), .C0(n8712), .Y(
        n8713) );
  AOI21X1TS U8844 ( .A0(n10147), .A1(n10397), .B0(n8713), .Y(n4548) );
  AOI31X1TS U8845 ( .A0(n9781), .A1(n9778), .A2(n11728), .B0(n12287), .Y(n8714) );
  OAI21X1TS U8846 ( .A0(n11722), .A1(n10250), .B0(n12543), .Y(n8715) );
  AOI32X1TS U8847 ( .A0(n11371), .A1(n8715), .A2(n9402), .B0(n11982), .B1(
        n8715), .Y(n8716) );
  AOI211X1TS U8848 ( .A0(n10237), .A1(n6655), .B0(n8714), .C0(n8716), .Y(n8717) );
  OAI2BB1X1TS U8849 ( .A0N(n12280), .A1N(n11760), .B0(n8717), .Y(n8718) );
  OAI32X1TS U8850 ( .A0(n8718), .A1(n10237), .A2(n9407), .B0(n12061), .B1(
        n8718), .Y(n8719) );
  OAI21X1TS U8851 ( .A0(n10969), .A1(n12433), .B0(n12298), .Y(n8720) );
  OAI211X1TS U8852 ( .A0(n10487), .A1(n11984), .B0(n8719), .C0(n8720), .Y(
        n5736) );
  AOI22X1TS U8853 ( .A0(n12180), .A1(n2535), .B0(n11953), .B1(n10680), .Y(
        n8721) );
  OAI211X1TS U8854 ( .A0(n10007), .A1(n1686), .B0(n1687), .C0(n8721), .Y(n8722) );
  OAI22X1TS U8855 ( .A0(n11637), .A1(n10695), .B0(n12565), .B1(n11643), .Y(
        n8723) );
  OAI211X1TS U8856 ( .A0(n10303), .A1(n2022), .B0(n1683), .C0(n1684), .Y(n8724) );
  AOI31X1TS U8857 ( .A0(n9764), .A1(n10689), .A2(n12563), .B0(n11949), .Y(
        n8725) );
  OAI22X1TS U8858 ( .A0(n10011), .A1(n1670), .B0(n1672), .B1(n10694), .Y(n8726) );
  AOI22X1TS U8859 ( .A0(n11955), .A1(n12186), .B0(n12192), .B1(n12646), .Y(
        n8727) );
  OAI211X1TS U8860 ( .A0(n10015), .A1(n1662), .B0(n1665), .C0(n8727), .Y(n8728) );
  NOR4XLTS U8861 ( .A(n1659), .B(n8725), .C(n8726), .D(n8728), .Y(n8729) );
  NAND3X1TS U8862 ( .A(n1654), .B(n8729), .C(n1655), .Y(n8730) );
  NOR4XLTS U8863 ( .A(n8722), .B(n8723), .C(n8724), .D(n8730), .Y(n1327) );
  OR4X1TS U8864 ( .A(n12344), .B(n12481), .C(n8180), .D(n9515), .Y(n8731) );
  OA22X1TS U8865 ( .A0(n8179), .A1(n10352), .B0(n8178), .B1(n11574), .Y(n8732)
         );
  OAI211X1TS U8866 ( .A0(n8175), .A1(n11575), .B0(n7978), .C0(n8732), .Y(n8733) );
  AOI211X1TS U8867 ( .A0(n10691), .A1(n8731), .B0(n8177), .C0(n8733), .Y(n8734) );
  NAND4X1TS U8868 ( .A(n7457), .B(n7269), .C(n8734), .D(n7596), .Y(n8735) );
  AOI22X1TS U8869 ( .A0(n8211), .A1(n12628), .B0(n8210), .B1(n10332), .Y(n8736) );
  AOI22X1TS U8870 ( .A0(n11133), .A1(n12178), .B0(n10102), .B1(n11945), .Y(
        n8737) );
  OAI211X1TS U8871 ( .A0(n8206), .A1(n12164), .B0(n8736), .C0(n8737), .Y(n8738) );
  NOR4XLTS U8872 ( .A(n8168), .B(n7575), .C(n8735), .D(n8738), .Y(n6932) );
  AOI2BB2X1TS U8873 ( .B0(n2914), .B1(n10264), .A0N(n9939), .A1N(n10207), .Y(
        n8739) );
  AOI2BB2X1TS U8874 ( .B0(n10527), .B1(n12140), .A0N(n12078), .A1N(n11888), 
        .Y(n8740) );
  OAI211X1TS U8875 ( .A0(sa21[6]), .A1(n8739), .B0(n2911), .C0(n8740), .Y(
        n8741) );
  AOI211X1TS U8876 ( .A0(n10263), .A1(n2319), .B0(n2906), .C0(n8741), .Y(n8742) );
  AOI32X1TS U8877 ( .A0(n9991), .A1(n8742), .A2(n12080), .B0(n11583), .B1(
        n8742), .Y(n8743) );
  AOI21X1TS U8878 ( .A0(n11847), .A1(n11100), .B0(n8743), .Y(n1695) );
  NOR3BX1TS U8879 ( .AN(n3322), .B(sa03[7]), .C(sa03[5]), .Y(n1987) );
  NAND3X1TS U8880 ( .A(n9066), .B(n9525), .C(n11816), .Y(n8744) );
  OAI2BB1X1TS U8881 ( .A0N(n11029), .A1N(n11828), .B0(n8744), .Y(n8745) );
  AOI21X1TS U8882 ( .A0(n11458), .A1(n10508), .B0(n11035), .Y(n8746) );
  AOI211X1TS U8883 ( .A0(n12452), .A1(n11827), .B0(n8746), .C0(n3027), .Y(
        n8747) );
  OAI21X1TS U8884 ( .A0(n12290), .A1(n10948), .B0(n10519), .Y(n8748) );
  NAND4BX1TS U8885 ( .AN(n3042), .B(n3065), .C(n8747), .D(n8748), .Y(n8749) );
  AOI211X1TS U8886 ( .A0(n11542), .A1(n3297), .B0(n8745), .C0(n8749), .Y(n2472) );
  AOI2BB2X1TS U8887 ( .B0(n12003), .B1(n12585), .A0N(n10393), .A1N(n11364), 
        .Y(n8750) );
  OAI211X1TS U8888 ( .A0(n4633), .A1(n10486), .B0(n8750), .C0(n4635), .Y(n8751) );
  OAI22X1TS U8889 ( .A0(n10837), .A1(n10910), .B0(n10393), .B1(n11411), .Y(
        n8752) );
  AOI211X1TS U8890 ( .A0(n10916), .A1(n4426), .B0(n4413), .C0(n8752), .Y(n8753) );
  AOI22X1TS U8891 ( .A0(n11231), .A1(n11739), .B0(n11743), .B1(n11357), .Y(
        n8754) );
  NAND4BX1TS U8892 ( .AN(n8751), .B(n8753), .C(n4421), .D(n8754), .Y(n3713) );
  OAI2BB2XLTS U8893 ( .B0(n11978), .B1(n6189), .A0N(n6046), .A1N(n10558), .Y(
        n8755) );
  AOI21X1TS U8894 ( .A0(n12575), .A1(n11676), .B0(n8755), .Y(n8756) );
  OAI21X1TS U8895 ( .A0(n10842), .A1(n9375), .B0(n10491), .Y(n8757) );
  OAI211X1TS U8896 ( .A0(n6039), .A1(n12495), .B0(n8756), .C0(n8757), .Y(n5814) );
  AOI31X1TS U8897 ( .A0(n9921), .A1(n12414), .A2(n9902), .B0(n12540), .Y(n8758) );
  OAI21X1TS U8898 ( .A0(n10813), .A1(n10133), .B0(n12620), .Y(n8759) );
  AOI32X1TS U8899 ( .A0(n9673), .A1(n8759), .A2(n12208), .B0(n12024), .B1(
        n8759), .Y(n8760) );
  OAI22X1TS U8900 ( .A0(n10769), .A1(n4492), .B0(n12206), .B1(n4856), .Y(n8761) );
  AOI22X1TS U8901 ( .A0(n11212), .A1(n10400), .B0(n4536), .B1(n10391), .Y(
        n8762) );
  OAI21X1TS U8902 ( .A0(n11767), .A1(n9118), .B0(n9691), .Y(n8763) );
  OAI211X1TS U8903 ( .A0(n10867), .A1(n12024), .B0(n8762), .C0(n8763), .Y(
        n8764) );
  OR4X1TS U8904 ( .A(n8758), .B(n8760), .C(n8761), .D(n8764), .Y(n3937) );
  AOI22X1TS U8905 ( .A0(n12331), .A1(n11513), .B0(n11519), .B1(n12151), .Y(
        n8765) );
  AOI211X1TS U8906 ( .A0(n12645), .A1(n2185), .B0(n2186), .C0(n2187), .Y(n8766) );
  AND4X1TS U8907 ( .A(n8765), .B(n2181), .C(n8766), .D(n2182), .Y(n8767) );
  AOI22X1TS U8908 ( .A0(n11003), .A1(n12186), .B0(n11507), .B1(n12195), .Y(
        n8768) );
  AOI22X1TS U8909 ( .A0(n9086), .A1(n1692), .B0(n11912), .B1(n2201), .Y(n8769)
         );
  OAI21X1TS U8910 ( .A0(n10607), .A1(n12556), .B0(n8769), .Y(n8770) );
  AOI211X1TS U8911 ( .A0(n12188), .A1(n11822), .B0(n2199), .C0(n8770), .Y(
        n8771) );
  AOI31X1TS U8912 ( .A0(sa32[6]), .A1(n2194), .A2(n1810), .B0(n2195), .Y(n8772) );
  NAND4X1TS U8913 ( .A(n8767), .B(n8768), .C(n8771), .D(n8772), .Y(n8773) );
  AOI22X1TS U8914 ( .A0(n1674), .A1(n2228), .B0(n12192), .B1(n1806), .Y(n8774)
         );
  AOI222XLTS U8915 ( .A0(n11919), .A1(n1802), .B0(n11051), .B1(n2213), .C0(
        n11501), .C1(n2224), .Y(n8775) );
  NAND4BX1TS U8916 ( .AN(n2226), .B(n8774), .C(n2227), .D(n8775), .Y(n8776) );
  NOR4XLTS U8917 ( .A(n1796), .B(n2178), .C(n8773), .D(n8776), .Y(n1374) );
  OAI22X1TS U8918 ( .A0(n11920), .A1(n10706), .B0(n11868), .B1(n10719), .Y(
        n8777) );
  AOI22X1TS U8919 ( .A0(n7491), .A1(n11139), .B0(n9542), .B1(n12632), .Y(n8778) );
  AOI31X1TS U8920 ( .A0(n9365), .A1(n9546), .A2(n11146), .B0(n7697), .Y(n8779)
         );
  OAI22X1TS U8921 ( .A0(n7690), .A1(n10343), .B0(n7667), .B1(n10338), .Y(n8780) );
  AOI211X1TS U8922 ( .A0(n7686), .A1(n10315), .B0(n7687), .C0(n8780), .Y(n8781) );
  OAI211X1TS U8923 ( .A0(n7681), .A1(n10066), .B0(n7683), .C0(n7684), .Y(n8782) );
  OAI21X1TS U8924 ( .A0(n11527), .A1(n10713), .B0(n7677), .Y(n8783) );
  NOR3X1TS U8925 ( .A(n7679), .B(n8782), .C(n8783), .Y(n8784) );
  NAND4X1TS U8926 ( .A(n8778), .B(n8779), .C(n8781), .D(n8784), .Y(n8785) );
  OAI22X1TS U8927 ( .A0(n7333), .A1(n9857), .B0(n9491), .B1(n11557), .Y(n8786)
         );
  NOR4XLTS U8928 ( .A(n7669), .B(n8777), .C(n8785), .D(n8786), .Y(n7306) );
  AOI22X1TS U8929 ( .A0(n12088), .A1(n10321), .B0(n7509), .B1(n10254), .Y(
        n8787) );
  AOI22X1TS U8930 ( .A0(n7765), .A1(n10017), .B0(n10622), .B1(n7128), .Y(n8788) );
  OAI211X1TS U8931 ( .A0(n10628), .A1(n9818), .B0(n8787), .C0(n8788), .Y(n8789) );
  AOI211X1TS U8932 ( .A0(n11564), .A1(n11444), .B0(n7529), .C0(n8789), .Y(
        n8790) );
  OAI22X1TS U8933 ( .A0(n11128), .A1(n10054), .B0(n12075), .B1(n12120), .Y(
        n8791) );
  OAI22X1TS U8934 ( .A0(n12321), .A1(n12335), .B0(n10033), .B1(n7536), .Y(
        n8792) );
  AOI22X1TS U8935 ( .A0(n10324), .A1(n10634), .B0(n11076), .B1(n12090), .Y(
        n8793) );
  OAI211X1TS U8936 ( .A0(n12306), .A1(n12319), .B0(n8793), .C0(n7870), .Y(
        n8794) );
  NOR4XLTS U8937 ( .A(n7865), .B(n8791), .C(n8792), .D(n8794), .Y(n8795) );
  OAI211X1TS U8938 ( .A0(n12102), .A1(n7520), .B0(n8790), .C0(n8795), .Y(n8796) );
  NOR4XLTS U8939 ( .A(n7742), .B(n7350), .C(n7861), .D(n8796), .Y(n6924) );
  OAI22X1TS U8940 ( .A0(n4656), .A1(n10815), .B0(n12396), .B1(n4120), .Y(n8797) );
  OAI22X1TS U8941 ( .A0(n11238), .A1(n4667), .B0(n10117), .B1(n4205), .Y(n8798) );
  OAI2BB2XLTS U8942 ( .B0(n4705), .B1(n10114), .A0N(n4698), .A1N(n11285), .Y(
        n8799) );
  OAI22X1TS U8943 ( .A0(n11993), .A1(n4087), .B0(n10113), .B1(n4121), .Y(n8800) );
  NOR4XLTS U8944 ( .A(n8797), .B(n8798), .C(n8799), .D(n8800), .Y(n8801) );
  OAI31X1TS U8945 ( .A0(sa22[2]), .A1(n9248), .A2(n12395), .B0(n4703), .Y(
        n8802) );
  OAI22X1TS U8946 ( .A0(n4204), .A1(n10811), .B0(n11400), .B1(n11296), .Y(
        n8803) );
  AOI211X1TS U8947 ( .A0(n12419), .A1(n12239), .B0(n8802), .C0(n8803), .Y(
        n8804) );
  AOI22X1TS U8948 ( .A0(n12229), .A1(n12236), .B0(n9638), .B1(n11309), .Y(
        n8805) );
  NAND4X1TS U8949 ( .A(n3877), .B(n8801), .C(n8804), .D(n8805), .Y(n8806) );
  OAI211X1TS U8950 ( .A0(n12429), .A1(n9110), .B0(n4208), .C0(n4209), .Y(n8807) );
  NOR4XLTS U8951 ( .A(n4429), .B(n4212), .C(n8806), .D(n8807), .Y(n3433) );
  OAI22X1TS U8952 ( .A0(n10469), .A1(n10923), .B0(n12424), .B1(n5920), .Y(
        n8808) );
  OAI22X1TS U8953 ( .A0(n11391), .A1(n6467), .B0(n10221), .B1(n6115), .Y(n8809) );
  OAI2BB2XLTS U8954 ( .B0(n6505), .B1(n10218), .A0N(n6498), .A1N(n11319), .Y(
        n8810) );
  OAI22X1TS U8955 ( .A0(n12040), .A1(n5887), .B0(n10217), .B1(n5921), .Y(n8811) );
  NOR4XLTS U8956 ( .A(n8808), .B(n8809), .C(n8810), .D(n8811), .Y(n8812) );
  OAI31X1TS U8957 ( .A0(n11201), .A1(n9444), .A2(n12423), .B0(n6503), .Y(n8813) );
  OAI22X1TS U8958 ( .A0(n6114), .A1(n10931), .B0(n11217), .B1(n11305), .Y(
        n8814) );
  AOI211X1TS U8959 ( .A0(n12407), .A1(n12250), .B0(n8813), .C0(n8814), .Y(
        n8815) );
  AOI22X1TS U8960 ( .A0(n12256), .A1(n12247), .B0(n9633), .B1(n11294), .Y(
        n8816) );
  NAND4X1TS U8961 ( .A(n5707), .B(n8812), .C(n8815), .D(n8816), .Y(n8817) );
  OAI211X1TS U8962 ( .A0(n12401), .A1(n9302), .B0(n6118), .C0(n6119), .Y(n8818) );
  NOR4XLTS U8963 ( .A(n6232), .B(n6122), .C(n8817), .D(n8818), .Y(n5230) );
  AOI22X1TS U8964 ( .A0(n9482), .A1(n11091), .B0(n11492), .B1(n9821), .Y(n8819) );
  AOI22X1TS U8965 ( .A0(n7964), .A1(n12470), .B0(n11086), .B1(n12636), .Y(
        n8820) );
  OAI211X1TS U8966 ( .A0(n12127), .A1(n7275), .B0(n8819), .C0(n8820), .Y(n8821) );
  AOI31X1TS U8967 ( .A0(sa02[0]), .A1(n9476), .A2(n12642), .B0(n8821), .Y(
        n8822) );
  NAND4X1TS U8968 ( .A(n7269), .B(n7268), .C(n7270), .D(n8822), .Y(n8823) );
  AOI22X1TS U8969 ( .A0(n12480), .A1(n7300), .B0(n9487), .B1(n10643), .Y(n8824) );
  AOI21X1TS U8970 ( .A0(n7296), .A1(n11504), .B0(n7297), .Y(n8825) );
  OAI31X1TS U8971 ( .A0(n12134), .A1(n9486), .A2(n12628), .B0(n11498), .Y(
        n8826) );
  NAND4X1TS U8972 ( .A(n7289), .B(n8824), .C(n8825), .D(n8826), .Y(n8827) );
  NOR4XLTS U8973 ( .A(n7264), .B(n7265), .C(n8823), .D(n8827), .Y(n1284) );
  AOI2BB2X1TS U8974 ( .B0(n10239), .B1(n2838), .A0N(n9935), .A1N(n10215), .Y(
        n8828) );
  AOI2BB2X1TS U8975 ( .B0(n10557), .B1(n12126), .A0N(n12086), .A1N(n11864), 
        .Y(n8829) );
  OAI211X1TS U8976 ( .A0(sa10[6]), .A1(n8828), .B0(n2835), .C0(n8829), .Y(
        n8830) );
  AOI211X1TS U8977 ( .A0(n11567), .A1(n10239), .B0(n2830), .C0(n8830), .Y(
        n8831) );
  AOI32X1TS U8978 ( .A0(n1926), .A1(n8831), .A2(n9980), .B0(n11571), .B1(n8831), .Y(n8832) );
  AOI21X1TS U8979 ( .A0(n1758), .A1(n11841), .B0(n8832), .Y(n1733) );
  NOR3BX1TS U8980 ( .AN(n5092), .B(n10308), .C(sa00[0]), .Y(n3673) );
  OAI2BB2XLTS U8981 ( .B0(n12039), .B1(n4386), .A0N(n4279), .A1N(n10374), .Y(
        n8833) );
  AOI21X1TS U8982 ( .A0(n12593), .A1(n11787), .B0(n8833), .Y(n8834) );
  OAI21X1TS U8983 ( .A0(n10928), .A1(n9179), .B0(n10433), .Y(n8835) );
  OAI211X1TS U8984 ( .A0(n4272), .A1(n12547), .B0(n8834), .C0(n8835), .Y(n3982) );
  NOR2X1TS U8985 ( .A(n12310), .B(n11011), .Y(n8836) );
  OAI22X1TS U8986 ( .A0(n2510), .A1(n10192), .B0(n8836), .B1(n11447), .Y(n8837) );
  AOI22X1TS U8987 ( .A0(n11560), .A1(n12451), .B0(n11441), .B1(n12623), .Y(
        n8838) );
  OAI211X1TS U8988 ( .A0(n10236), .A1(n12117), .B0(n2766), .C0(n8838), .Y(
        n8839) );
  OAI22X1TS U8989 ( .A0(n11036), .A1(n11857), .B0(n11835), .B1(n11448), .Y(
        n8840) );
  AOI21X1TS U8990 ( .A0(n12106), .A1(n11815), .B0(n2160), .Y(n8841) );
  OAI31X1TS U8991 ( .A0(n3315), .A1(n11460), .A2(sa03[7]), .B0(n8841), .Y(
        n8842) );
  NOR4XLTS U8992 ( .A(n8837), .B(n8839), .C(n8840), .D(n8842), .Y(n2044) );
  AOI22X1TS U8993 ( .A0(n10538), .A1(n12598), .B0(n10272), .B1(n11490), .Y(
        n8843) );
  OAI21X1TS U8994 ( .A0(n11935), .A1(n11153), .B0(n9984), .Y(n8844) );
  NAND4X1TS U8995 ( .A(n2340), .B(n1840), .C(n8843), .D(n8844), .Y(n8845) );
  AOI211X1TS U8996 ( .A0(n10300), .A1(n12372), .B0(n2309), .C0(n8845), .Y(
        n2395) );
  AOI22X1TS U8997 ( .A0(n11678), .A1(n10953), .B0(n11675), .B1(n10145), .Y(
        n8846) );
  AOI31X1TS U8998 ( .A0(n10820), .A1(n5315), .A2(n12198), .B0(n11689), .Y(
        n8847) );
  AOI211X1TS U8999 ( .A0(n6699), .A1(n11336), .B0(n6175), .C0(n8847), .Y(n8848) );
  OAI211X1TS U9000 ( .A0(n10980), .A1(n6043), .B0(n8846), .C0(n8848), .Y(n8849) );
  AOI22X1TS U9001 ( .A0(n10496), .A1(n9969), .B0(n11207), .B1(n5418), .Y(n8850) );
  OAI21X1TS U9002 ( .A0(n11377), .A1(n10559), .B0(n11979), .Y(n8851) );
  NAND4X1TS U9003 ( .A(n6163), .B(n5634), .C(n8850), .D(n8851), .Y(n8852) );
  OAI22X1TS U9004 ( .A0(n5413), .A1(n10989), .B0(n10500), .B1(n5414), .Y(n8853) );
  AOI211X1TS U9005 ( .A0(n11697), .A1(n12449), .B0(n6578), .C0(n8853), .Y(
        n8854) );
  OAI211X1TS U9006 ( .A0(n5310), .A1(n10154), .B0(n6144), .C0(n8854), .Y(n8855) );
  NOR4XLTS U9007 ( .A(n5280), .B(n8849), .C(n8852), .D(n8855), .Y(n5238) );
  AOI22X1TS U9008 ( .A0(n11703), .A1(n10401), .B0(n10459), .B1(n10798), .Y(
        n8856) );
  AOI31X1TS U9009 ( .A0(n11382), .A1(n3647), .A2(n12541), .B0(n11756), .Y(
        n8857) );
  AOI211X1TS U9010 ( .A0(n4837), .A1(n3969), .B0(n4561), .C0(n8857), .Y(n8858)
         );
  OAI211X1TS U9011 ( .A0(n11714), .A1(n4509), .B0(n8856), .C0(n8858), .Y(n8859) );
  AOI22X1TS U9012 ( .A0(n3640), .A1(n10134), .B0(n10876), .B1(n3918), .Y(n8860) );
  OAI21X1TS U9013 ( .A0(n10138), .A1(n9691), .B0(n11374), .Y(n8861) );
  NAND4X1TS U9014 ( .A(n4548), .B(n3961), .C(n8860), .D(n8861), .Y(n8862) );
  OAI22X1TS U9015 ( .A0(n3913), .A1(n10861), .B0(n12571), .B1(n3914), .Y(n8863) );
  AOI211X1TS U9016 ( .A0(n12202), .A1(n11767), .B0(n4824), .C0(n8863), .Y(
        n8864) );
  OAI211X1TS U9017 ( .A0(n9677), .A1(n12380), .B0(n4526), .C0(n8864), .Y(n8865) );
  NOR4XLTS U9018 ( .A(n3637), .B(n8859), .C(n8862), .D(n8865), .Y(n3390) );
  NOR3X1TS U9019 ( .A(sa21[2]), .B(n9068), .C(n11907), .Y(n8866) );
  AOI211X1TS U9020 ( .A0(n12139), .A1(n11136), .B0(n2390), .C0(n8866), .Y(
        n8867) );
  OAI22X1TS U9021 ( .A0(n11900), .A1(n11888), .B0(n2311), .B1(n11905), .Y(
        n8868) );
  OAI22X1TS U9022 ( .A0(n10547), .A1(n2932), .B0(n10211), .B1(n2392), .Y(n8869) );
  OAI22X1TS U9023 ( .A0(n2881), .A1(n10978), .B0(n2920), .B1(n12485), .Y(n8870) );
  OAI22X1TS U9024 ( .A0(n11435), .A1(n9113), .B0(n2313), .B1(n10977), .Y(n8871) );
  NOR4XLTS U9025 ( .A(n8868), .B(n8869), .C(n8870), .D(n8871), .Y(n8872) );
  NAND4X1TS U9026 ( .A(n2080), .B(n2393), .C(n8867), .D(n8872), .Y(n8873) );
  OAI22X1TS U9027 ( .A0(n11482), .A1(n2346), .B0(n2379), .B1(n12475), .Y(n8874) );
  AOI211X1TS U9028 ( .A0(n12146), .A1(n10284), .B0(n2304), .C0(n8874), .Y(
        n8875) );
  AOI32X1TS U9029 ( .A0(n12482), .A1(n8875), .A2(n12176), .B0(n10649), .B1(
        n8875), .Y(n8876) );
  NOR4XLTS U9030 ( .A(n2672), .B(n2402), .C(n8873), .D(n8876), .Y(n1470) );
  AOI31X1TS U9031 ( .A0(n10426), .A1(n9659), .A2(n3871), .B0(n10843), .Y(n8877) );
  AOI32X1TS U9032 ( .A0(n3866), .A1(n3865), .A2(n3864), .B0(n11345), .B1(n3865), .Y(n8878) );
  AOI22X1TS U9033 ( .A0(n3555), .A1(n11332), .B0(n12221), .B1(n12515), .Y(
        n8879) );
  AOI22X1TS U9034 ( .A0(n10832), .A1(n12262), .B0(n3862), .B1(n10915), .Y(
        n8880) );
  NAND4X1TS U9035 ( .A(n3861), .B(n3859), .C(n8879), .D(n8880), .Y(n8881) );
  AOI211X1TS U9036 ( .A0(n11332), .A1(n10906), .B0(n3856), .C0(n8881), .Y(
        n8882) );
  NAND4X1TS U9037 ( .A(n3854), .B(n3853), .C(n8882), .D(n3852), .Y(n8883) );
  NOR2X1TS U9038 ( .A(n12059), .B(n12222), .Y(n8884) );
  OAI22X1TS U9039 ( .A0(n3868), .A1(n11262), .B0(n8884), .B1(n10838), .Y(n8885) );
  NOR4XLTS U9040 ( .A(n8877), .B(n8878), .C(n8883), .D(n8885), .Y(n3338) );
  XOR2X1TS U9041 ( .A(n1781), .B(n1548), .Y(n3429) );
  XOR2X1TS U9042 ( .A(n1648), .B(n1533), .Y(n5226) );
  XOR2X1TS U9043 ( .A(n1486), .B(n1417), .Y(n1323) );
  OAI22X1TS U9044 ( .A0(n12011), .A1(n5674), .B0(n6341), .B1(n11736), .Y(n8886) );
  AOI2BB2X1TS U9045 ( .B0(n11354), .B1(n5670), .A0N(n5668), .A1N(n12286), .Y(
        n8887) );
  OAI21X1TS U9046 ( .A0(n5676), .A1(n11735), .B0(n8887), .Y(n8888) );
  AOI211X1TS U9047 ( .A0(n10968), .A1(n5677), .B0(n8886), .C0(n8888), .Y(n8889) );
  NAND4X1TS U9048 ( .A(n5660), .B(n11730), .C(n12004), .D(n5662), .Y(n8890) );
  AOI222XLTS U9049 ( .A0(n11347), .A1(n9973), .B0(n10970), .B1(n9978), .C0(
        n10194), .C1(n10963), .Y(n8891) );
  NAND4BX1TS U9050 ( .AN(n5648), .B(n5652), .C(n8891), .D(n5650), .Y(n8892) );
  AOI211X1TS U9051 ( .A0(n10946), .A1(n8890), .B0(n5643), .C0(n8892), .Y(n8893) );
  NAND4X1TS U9052 ( .A(n8889), .B(n5664), .C(n8893), .D(n5644), .Y(n1777) );
  OAI21X1TS U9053 ( .A0(n10098), .A1(n11952), .B0(n7993), .Y(n8894) );
  OAI31X1TS U9054 ( .A0(n8364), .A1(n9593), .A2(n10352), .B0(n7627), .Y(n8895)
         );
  AOI211X1TS U9055 ( .A0(n10642), .A1(n12479), .B0(n8894), .C0(n8895), .Y(
        n8896) );
  NOR2X1TS U9056 ( .A(n10101), .B(n10090), .Y(n8897) );
  OAI22X1TS U9057 ( .A0(n11640), .A1(n8897), .B0(n10085), .B1(n8206), .Y(n8898) );
  AOI211X1TS U9058 ( .A0(n11579), .A1(n7296), .B0(n7576), .C0(n8898), .Y(n8899) );
  AOI22X1TS U9059 ( .A0(n7455), .A1(n7979), .B0(n11133), .B1(n7467), .Y(n8900)
         );
  OAI211X1TS U9060 ( .A0(n8190), .A1(n11178), .B0(n8259), .C0(n8900), .Y(n8901) );
  OAI21X1TS U9061 ( .A0(n11493), .A1(n10306), .B0(n12473), .Y(n8902) );
  OAI211X1TS U9062 ( .A0(n7974), .A1(n8231), .B0(n8358), .C0(n8902), .Y(n8903)
         );
  AOI211X1TS U9063 ( .A0(n12177), .A1(n10311), .B0(n8901), .C0(n8903), .Y(
        n8904) );
  NAND4X1TS U9064 ( .A(n7616), .B(n8896), .C(n8899), .D(n8904), .Y(n8905) );
  AOI22X1TS U9065 ( .A0(n8203), .A1(n8240), .B0(n10301), .B1(n8370), .Y(n8906)
         );
  NAND3X1TS U9066 ( .A(n7617), .B(n7270), .C(n8906), .Y(n8907) );
  NOR4XLTS U9067 ( .A(n8168), .B(n7265), .C(n8905), .D(n8907), .Y(n1273) );
  OAI22X1TS U9068 ( .A0(n11101), .A1(n10065), .B0(n10719), .B1(n9858), .Y(
        n8908) );
  AOI211X1TS U9069 ( .A0(n12633), .A1(n11855), .B0(n8301), .C0(n8908), .Y(
        n8909) );
  NAND3X1TS U9070 ( .A(n11150), .B(n10341), .C(n10077), .Y(n8910) );
  OAI211X1TS U9071 ( .A0(n7331), .A1(n10648), .B0(n8909), .C0(n8910), .Y(n8911) );
  OAI22X1TS U9072 ( .A0(n11867), .A1(n7681), .B0(n10338), .B1(n8306), .Y(n8912) );
  OAI22X1TS U9073 ( .A0(n11521), .A1(n7729), .B0(n11511), .B1(n7834), .Y(n8913) );
  NOR2X1TS U9074 ( .A(n11097), .B(n11553), .Y(n8914) );
  AOI22X1TS U9075 ( .A0(n10282), .A1(n7838), .B0(n7836), .B1(n11896), .Y(n8915) );
  OAI211X1TS U9076 ( .A0(n11559), .A1(n8914), .B0(n8915), .C0(n8034), .Y(n8916) );
  AOI211X1TS U9077 ( .A0(n11928), .A1(n8286), .B0(n8913), .C0(n8916), .Y(n8917) );
  OAI22X1TS U9078 ( .A0(n11509), .A1(n11108), .B0(n11903), .B1(n10029), .Y(
        n8918) );
  NOR3X1TS U9079 ( .A(n7669), .B(n7653), .C(n8918), .Y(n8919) );
  NAND4X1TS U9080 ( .A(n8917), .B(n7319), .C(n7307), .D(n8919), .Y(n8920) );
  NOR4XLTS U9081 ( .A(n7811), .B(n7646), .C(n8912), .D(n8920), .Y(n8921) );
  NAND2X1TS U9082 ( .A(n7683), .B(n8921), .Y(n8922) );
  AOI211X1TS U9083 ( .A0(n10081), .A1(n11592), .B0(n8911), .C0(n8922), .Y(
        n1515) );
  OAI22X1TS U9084 ( .A0(n7246), .A1(n12559), .B0(n10678), .B1(n9805), .Y(n8923) );
  AO22X1TS U9085 ( .A0(n7570), .A1(n11564), .B0(n7128), .B1(n11569), .Y(n8924)
         );
  OAI211X1TS U9086 ( .A0(n7365), .A1(n11044), .B0(n7567), .C0(n7370), .Y(n8925) );
  AOI21X1TS U9087 ( .A0(n7564), .A1(n10634), .B0(n8925), .Y(n8926) );
  OAI22X1TS U9088 ( .A0(n12083), .A1(n11807), .B0(n11114), .B1(n11801), .Y(
        n8927) );
  OAI211X1TS U9089 ( .A0(n10683), .A1(n11872), .B0(n7561), .C0(n7562), .Y(
        n8928) );
  OAI31X1TS U9090 ( .A0(n7512), .A1(n9842), .A2(sa13[2]), .B0(n7563), .Y(n8929) );
  NOR4XLTS U9091 ( .A(n7556), .B(n8927), .C(n8928), .D(n8929), .Y(n8930) );
  OAI211X1TS U9092 ( .A0(n7252), .A1(n12103), .B0(n8926), .C0(n8930), .Y(n8931) );
  NOR3X1TS U9093 ( .A(n8923), .B(n8924), .C(n8931), .Y(n8932) );
  NAND4X1TS U9094 ( .A(n7223), .B(n7502), .C(n8932), .D(n7112), .Y(n1597) );
  NOR3BX1TS U9095 ( .AN(n6719), .B(sa30[5]), .C(n10716), .Y(n5297) );
  NOR3BX1TS U9096 ( .AN(n3191), .B(sa21[7]), .C(n10064), .Y(n1845) );
  NAND2BX1TS U9097 ( .AN(n9070), .B(n9066), .Y(n11021) );
  AOI2BB2X1TS U9098 ( .B0(n12050), .B1(n5931), .A0N(n10541), .A1N(n11289), .Y(
        n8933) );
  OAI211X1TS U9099 ( .A0(n6505), .A1(n10449), .B0(n8933), .C0(n6507), .Y(n8934) );
  OAI22X1TS U9100 ( .A0(n10929), .A1(n10873), .B0(n10541), .B1(n11216), .Y(
        n8935) );
  AOI211X1TS U9101 ( .A0(n10869), .A1(n6269), .B0(n6256), .C0(n8935), .Y(n8936) );
  AOI22X1TS U9102 ( .A0(n11414), .A1(n11712), .B0(n11704), .B1(n11294), .Y(
        n8937) );
  NAND4BX1TS U9103 ( .AN(n8934), .B(n8936), .C(n6264), .D(n8937), .Y(n5534) );
  AOI32X1TS U9104 ( .A0(n9662), .A1(n3764), .A2(n9111), .B0(n10816), .B1(n3764), .Y(n8938) );
  AOI211X1TS U9105 ( .A0(n11731), .A1(n12231), .B0(n3765), .C0(n8938), .Y(
        n8939) );
  OAI22X1TS U9106 ( .A0(n10131), .A1(n3768), .B0(n3591), .B1(n11316), .Y(n8940) );
  OAI22X1TS U9107 ( .A0(n10810), .A1(n3773), .B0(n11302), .B1(n11298), .Y(
        n8941) );
  AOI22X1TS U9108 ( .A0(n12507), .A1(n11733), .B0(n11394), .B1(n12579), .Y(
        n8942) );
  AOI21X1TS U9109 ( .A0(n10438), .A1(n10823), .B0(n12398), .Y(n8943) );
  AOI211X1TS U9110 ( .A0(n11322), .A1(n10828), .B0(n8943), .C0(n3754), .Y(
        n8944) );
  OAI31X1TS U9111 ( .A0(n10443), .A1(n12245), .A2(n12229), .B0(n12238), .Y(
        n8945) );
  NAND4X1TS U9112 ( .A(n3747), .B(n8942), .C(n8944), .D(n8945), .Y(n8946) );
  NOR4BX1TS U9113 ( .AN(n8939), .B(n8940), .C(n8941), .D(n8946), .Y(n8947) );
  AND4X1TS U9114 ( .A(n3564), .B(n8947), .C(n3741), .D(n3740), .Y(n1595) );
  AOI32X1TS U9115 ( .A0(n9667), .A1(n3698), .A2(n9103), .B0(n10845), .B1(n3698), .Y(n8948) );
  AOI211X1TS U9116 ( .A0(n11749), .A1(n12254), .B0(n3699), .C0(n8948), .Y(
        n8949) );
  OAI22X1TS U9117 ( .A0(n10139), .A1(n3702), .B0(n3552), .B1(n11364), .Y(n8950) );
  OAI22X1TS U9118 ( .A0(n10837), .A1(n3707), .B0(n11351), .B1(n11344), .Y(
        n8951) );
  AOI22X1TS U9119 ( .A0(n12522), .A1(n11751), .B0(n11406), .B1(n12587), .Y(
        n8952) );
  AOI21X1TS U9120 ( .A0(n10446), .A1(n10850), .B0(n12406), .Y(n8953) );
  AOI211X1TS U9121 ( .A0(n11370), .A1(n10856), .B0(n8953), .C0(n3688), .Y(
        n8954) );
  OAI31X1TS U9122 ( .A0(n10450), .A1(n12267), .A2(n12253), .B0(n12261), .Y(
        n8955) );
  NAND4X1TS U9123 ( .A(n3681), .B(n8952), .C(n8954), .D(n8955), .Y(n8956) );
  NOR4BX1TS U9124 ( .AN(n8949), .B(n8950), .C(n8951), .D(n8956), .Y(n8957) );
  AND4X1TS U9125 ( .A(n3525), .B(n8957), .C(n3675), .D(n3674), .Y(n1637) );
  NAND2BX1TS U9126 ( .AN(n4783), .B(n4281), .Y(n4245) );
  NOR3BX1TS U9127 ( .AN(n4920), .B(n9896), .C(n10752), .Y(n3499) );
  NOR3BX1TS U9128 ( .AN(n3251), .B(n10323), .C(sa10[5]), .Y(n1908) );
  NAND2X1TS U9129 ( .A(n10329), .B(n11873), .Y(n8958) );
  AOI22X1TS U9130 ( .A0(n7757), .A1(n12313), .B0(n11455), .B1(n8958), .Y(n8959) );
  OAI22X1TS U9131 ( .A0(n7755), .A1(n12084), .B0(n9829), .B1(n12322), .Y(n8960) );
  AOI22X1TS U9132 ( .A0(n11450), .A1(n11077), .B0(n7753), .B1(n10632), .Y(
        n8961) );
  OAI211X1TS U9133 ( .A0(n12304), .A1(n10627), .B0(n7561), .C0(n8961), .Y(
        n8962) );
  OAI211X1TS U9134 ( .A0(n12559), .A1(n10608), .B0(n7754), .C0(n7104), .Y(
        n8963) );
  NOR4XLTS U9135 ( .A(n7533), .B(n8960), .C(n8962), .D(n8963), .Y(n8964) );
  NAND4X1TS U9136 ( .A(n7354), .B(n7746), .C(n8959), .D(n8964), .Y(n8965) );
  OAI31X1TS U9137 ( .A0(n11037), .A1(n11564), .A2(n12638), .B0(n12314), .Y(
        n8966) );
  OAI211X1TS U9138 ( .A0(n7770), .A1(n10005), .B0(n7771), .C0(n8966), .Y(n8967) );
  NOR4XLTS U9139 ( .A(n7742), .B(n7743), .C(n8965), .D(n8967), .Y(n6925) );
  XOR2X1TS U9140 ( .A(n6935), .B(n1645), .Y(n6986) );
  XOR2X1TS U9141 ( .A(n6984), .B(n9155), .Y(n6936) );
  XOR2X1TS U9142 ( .A(n1407), .B(n1401), .Y(n1472) );
  XOR2X1TS U9143 ( .A(n6933), .B(n1566), .Y(n6942) );
  XOR2X1TS U9144 ( .A(n5159), .B(n1773), .Y(n5213) );
  XOR2X1TS U9145 ( .A(n3433), .B(n9084), .Y(n3384) );
  XOR2X1TS U9146 ( .A(n5230), .B(n9271), .Y(n5180) );
  XOR2X1TS U9147 ( .A(n3372), .B(n1784), .Y(n3422) );
  XOR2X1TS U9148 ( .A(n5166), .B(n1770), .Y(n5219) );
  OAI22X1TS U9149 ( .A0(n10771), .A1(n3962), .B0(n11381), .B1(n10407), .Y(
        n8968) );
  OAI22X1TS U9150 ( .A0(n3962), .A1(n12572), .B0(n3963), .B1(n10775), .Y(n8969) );
  OAI211X1TS U9151 ( .A0(n12413), .A1(n10777), .B0(n3960), .C0(n3961), .Y(
        n8970) );
  AOI211X1TS U9152 ( .A0(n12032), .A1(n3927), .B0(n8969), .C0(n8970), .Y(n8971) );
  OAI22X1TS U9153 ( .A0(n9670), .A1(n12024), .B0(n12567), .B1(n12382), .Y(
        n8972) );
  OAI22X1TS U9154 ( .A0(n10782), .A1(n3967), .B0(n3916), .B1(n12571), .Y(n8973) );
  AOI211X1TS U9155 ( .A0(n12029), .A1(n11249), .B0(n8972), .C0(n8973), .Y(
        n8974) );
  NAND4X1TS U9156 ( .A(n3632), .B(n8971), .C(n3966), .D(n8974), .Y(n8975) );
  NOR4XLTS U9157 ( .A(n3938), .B(n3937), .C(n8968), .D(n8975), .Y(n1993) );
  OAI22X1TS U9158 ( .A0(n10603), .A1(n10304), .B0(n2014), .B1(n11045), .Y(
        n8976) );
  OAI22X1TS U9159 ( .A0(n2014), .A1(n9968), .B0(n2012), .B1(n12554), .Y(n8977)
         );
  AOI211X1TS U9160 ( .A0(n9748), .A1(n12181), .B0(n2010), .C0(n8977), .Y(n8978) );
  NAND4X1TS U9161 ( .A(n2008), .B(n1799), .C(n8978), .D(n2006), .Y(n8979) );
  AOI22X1TS U9162 ( .A0(n10610), .A1(n2023), .B0(n1802), .B1(n12153), .Y(n8980) );
  AOI22X1TS U9163 ( .A0(n12182), .A1(n11594), .B0(n11157), .B1(n12187), .Y(
        n8981) );
  AOI22X1TS U9164 ( .A0(n1671), .A1(n11056), .B0(n11919), .B1(n12324), .Y(
        n8982) );
  NAND4X1TS U9165 ( .A(n8980), .B(n1684), .C(n8981), .D(n8982), .Y(n8983) );
  NOR4XLTS U9166 ( .A(n2002), .B(n8976), .C(n8979), .D(n8983), .Y(n1355) );
  AOI22X1TS U9167 ( .A0(n5617), .A1(n11336), .B0(n11980), .B1(n10951), .Y(
        n8984) );
  OAI22X1TS U9168 ( .A0(n11673), .A1(n9942), .B0(n5291), .B1(n6010), .Y(n8985)
         );
  AOI211X1TS U9169 ( .A0(n9953), .A1(n11669), .B0(n5611), .C0(n8985), .Y(n8986) );
  CLKINVX1TS U9170 ( .A(n5416), .Y(n8987) );
  AOI22X1TS U9171 ( .A0(n5614), .A1(n10141), .B0(n11229), .B1(n8987), .Y(n8988) );
  NAND4X1TS U9172 ( .A(n8984), .B(n5277), .C(n8986), .D(n8988), .Y(n8989) );
  OAI22X1TS U9173 ( .A0(n5641), .A1(n5424), .B0(n5639), .B1(n10189), .Y(n8990)
         );
  AOI211X1TS U9174 ( .A0(n10842), .A1(n9970), .B0(n5637), .C0(n8990), .Y(n8991) );
  OAI211X1TS U9175 ( .A0(n9288), .A1(n9941), .B0(n5634), .C0(n8991), .Y(n8992)
         );
  NOR4XLTS U9176 ( .A(n5604), .B(n5605), .C(n8989), .D(n8992), .Y(n1536) );
  AOI22X1TS U9177 ( .A0(n3822), .A1(n11273), .B0(n11810), .B1(n10799), .Y(
        n8993) );
  OAI22X1TS U9178 ( .A0(n11387), .A1(n9920), .B0(n3493), .B1(n4243), .Y(n8994)
         );
  AOI211X1TS U9179 ( .A0(n9904), .A1(n12045), .B0(n3816), .C0(n8994), .Y(n8995) );
  CLKINVX1TS U9180 ( .A(n3618), .Y(n8996) );
  AOI22X1TS U9181 ( .A0(n3819), .A1(n10159), .B0(n10883), .B1(n8996), .Y(n8997) );
  NAND4X1TS U9182 ( .A(n8993), .B(n3479), .C(n8995), .D(n8997), .Y(n8998) );
  OAI22X1TS U9183 ( .A0(n3846), .A1(n10789), .B0(n3844), .B1(n10120), .Y(n8999) );
  AOI211X1TS U9184 ( .A0(n10927), .A1(n9918), .B0(n3842), .C0(n8999), .Y(n9000) );
  OAI211X1TS U9185 ( .A0(n3628), .A1(n9919), .B0(n3839), .C0(n9000), .Y(n9001)
         );
  NOR4XLTS U9186 ( .A(n3809), .B(n3810), .C(n8998), .D(n9001), .Y(n1551) );
  CLKINVX1TS U9187 ( .A(n2058), .Y(n9002) );
  AOI22X1TS U9188 ( .A0(n9094), .A1(n10228), .B0(n2055), .B1(n11543), .Y(n9003) );
  OAI211X1TS U9189 ( .A0(n11548), .A1(n9002), .B0(n2053), .C0(n9003), .Y(n9004) );
  OAI22X1TS U9190 ( .A0(n2060), .A1(n11853), .B0(n2059), .B1(n12099), .Y(n9005) );
  NOR4XLTS U9191 ( .A(n2047), .B(n2048), .C(n9004), .D(n9005), .Y(n9006) );
  AOI22X1TS U9192 ( .A0(n10224), .A1(n9955), .B0(n2070), .B1(n11041), .Y(n9007) );
  NAND4X1TS U9193 ( .A(n11554), .B(n2073), .C(n11859), .D(n2074), .Y(n9008) );
  AOI22X1TS U9194 ( .A0(n9091), .A1(n9008), .B0(n11042), .B1(n11542), .Y(n9009) );
  OAI211X1TS U9195 ( .A0(n12315), .A1(n10598), .B0(n9007), .C0(n9009), .Y(
        n9010) );
  NOR3X1TS U9196 ( .A(n2043), .B(n2063), .C(n9010), .Y(n9011) );
  NAND3X1TS U9197 ( .A(n2044), .B(n9006), .C(n9011), .Y(n1331) );
  NAND2BX1TS U9198 ( .AN(n12654), .B(n11969), .Y(n1259) );
  OAI31X1TS U9199 ( .A0(n10068), .A1(n7630), .A2(n12155), .B0(n7631), .Y(n9012) );
  OAI21X1TS U9200 ( .A0(n10702), .A1(n7460), .B0(n9822), .Y(n9013) );
  OAI211X1TS U9201 ( .A0(n7960), .A1(n11586), .B0(n7627), .C0(n9013), .Y(n9014) );
  AOI211X1TS U9202 ( .A0(n11580), .A1(n12625), .B0(n9012), .C0(n9014), .Y(
        n9015) );
  AOI22X1TS U9203 ( .A0(n11497), .A1(n7594), .B0(n7593), .B1(n12343), .Y(n9016) );
  AOI21X1TS U9204 ( .A0(n8209), .A1(n12165), .B0(n12170), .Y(n9017) );
  OAI22X1TS U9205 ( .A0(n7587), .A1(n9527), .B0(n7585), .B1(n12158), .Y(n9018)
         );
  AOI211X1TS U9206 ( .A0(n7582), .A1(n12626), .B0(n9017), .C0(n9018), .Y(n9019) );
  AOI22X1TS U9207 ( .A0(n7447), .A1(n9481), .B0(n11093), .B1(n12641), .Y(n9020) );
  NAND4X1TS U9208 ( .A(n9016), .B(n7578), .C(n9019), .D(n9020), .Y(n9021) );
  NOR4XLTS U9209 ( .A(n7575), .B(n7264), .C(n7576), .D(n9021), .Y(n9022) );
  NAND3X1TS U9210 ( .A(n9015), .B(n7574), .C(n9022), .Y(n9023) );
  AOI211X1TS U9211 ( .A0(n10302), .A1(n9486), .B0(n7632), .C0(n9023), .Y(n1305) );
  AOI211X1TS U9212 ( .A0(n9761), .A1(n11111), .B0(n2089), .C0(n2088), .Y(n9024) );
  AOI32X1TS U9213 ( .A0(n10672), .A1(n9024), .A2(n1716), .B0(n12483), .B1(
        n9024), .Y(n9025) );
  AOI211X1TS U9214 ( .A0(n11104), .A1(n12600), .B0(n2083), .C0(n9025), .Y(
        n9026) );
  NAND4X1TS U9215 ( .A(n2081), .B(n2079), .C(n2080), .D(n9026), .Y(n9027) );
  AOI211X1TS U9216 ( .A0(n2898), .A1(n10727), .B0(n12137), .C0(n2100), .Y(
        n9028) );
  NAND2X1TS U9217 ( .A(n11141), .B(n10276), .Y(n9029) );
  AOI22X1TS U9218 ( .A0(n9729), .A1(n9029), .B0(n2096), .B1(n11847), .Y(n9030)
         );
  AOI22X1TS U9219 ( .A0(n11110), .A1(n2093), .B0(n11937), .B1(n2094), .Y(n9031) );
  OAI211X1TS U9220 ( .A0(n11889), .A1(n9028), .B0(n9030), .C0(n9031), .Y(n9032) );
  NOR4XLTS U9221 ( .A(n2075), .B(n2076), .C(n9027), .D(n9032), .Y(n1424) );
  XOR2X1TS U9222 ( .A(n9553), .B(text_in_r[3]), .Y(n9033) );
  AOI22X1TS U9223 ( .A0(n1455), .A1(n9083), .B0(n1454), .B1(n2229), .Y(n9034)
         );
  XOR2X1TS U9224 ( .A(n9034), .B(n1375), .Y(n9035) );
  XOR2X1TS U9225 ( .A(n9553), .B(n1352), .Y(n9036) );
  XOR2X1TS U9226 ( .A(n9035), .B(n9036), .Y(n9037) );
  OAI22X1TS U9227 ( .A0(n9033), .A1(n12690), .B0(n12753), .B1(n9037), .Y(N35)
         );
  INVXLTS U9228 ( .A(n9038), .Y(n9039) );
  INVXLTS U9229 ( .A(n1198), .Y(n9040) );
  INVXLTS U9230 ( .A(n9040), .Y(n9041) );
  INVX1TS U9231 ( .A(n3345), .Y(n9077) );
  INVX1TS U9232 ( .A(n5217), .Y(n12658) );
  INVX1TS U9233 ( .A(n5147), .Y(n9268) );
  INVX2TS U9234 ( .A(n1294), .Y(n9784) );
  CLKINVX2TS U9235 ( .A(n1456), .Y(n9772) );
  INVXLTS U9236 ( .A(n6980), .Y(n9128) );
  INVXLTS U9237 ( .A(n5182), .Y(n9210) );
  INVXLTS U9238 ( .A(n3386), .Y(n9195) );
  INVX2TS U9239 ( .A(n1615), .Y(n9768) );
  INVX2TS U9240 ( .A(n1540), .Y(n9202) );
  CLKINVX1TS U9241 ( .A(n1529), .Y(n9213) );
  INVXLTS U9242 ( .A(n3346), .Y(n9188) );
  INVXLTS U9243 ( .A(n5186), .Y(n9117) );
  CLKINVX1TS U9244 ( .A(n3330), .Y(n9131) );
  CLKINVX2TS U9245 ( .A(n5233), .Y(n9280) );
  CLKINVX1TS U9246 ( .A(n3441), .Y(n9185) );
  INVXLTS U9247 ( .A(n5140), .Y(n9207) );
  CLKINVX2TS U9248 ( .A(n3436), .Y(n9093) );
  CLKINVX1TS U9249 ( .A(n1581), .Y(n9171) );
  AOI22X1TS U9250 ( .A0(n12647), .A1(n9086), .B0(n10610), .B1(n9748), .Y(n2219) );
  AOI211X1TS U9251 ( .A0(n11395), .A1(n12449), .B0(n5292), .C0(n6007), .Y(
        n6005) );
  AOI211X1TS U9252 ( .A0(n11677), .A1(n12448), .B0(n5611), .C0(n6036), .Y(
        n6034) );
  AOI211X1TS U9253 ( .A0(n11218), .A1(n12376), .B0(n3494), .C0(n4240), .Y(
        n4238) );
  INVX1TS U9254 ( .A(n8175), .Y(n9510) );
  CLKINVX1TS U9255 ( .A(n12031), .Y(n10455) );
  INVX1TS U9256 ( .A(n7734), .Y(n10723) );
  CLKINVX1TS U9257 ( .A(n4020), .Y(n9122) );
  CLKINVX2TS U9258 ( .A(n12032), .Y(n10456) );
  AOI22X1TS U9259 ( .A0(n12199), .A1(n10875), .B0(n11779), .B1(n11374), .Y(
        n5097) );
  CLKINVX2TS U9260 ( .A(n7163), .Y(n11820) );
  CLKINVX2TS U9261 ( .A(n3583), .Y(n12429) );
  CLKINVX1TS U9262 ( .A(n5381), .Y(n12402) );
  AOI22X1TS U9263 ( .A0(n12528), .A1(n12271), .B0(n11317), .B1(n5392), .Y(
        n5713) );
  INVX2TS U9264 ( .A(n10817), .Y(n10772) );
  CLKINVX2TS U9265 ( .A(n1938), .Y(n12347) );
  CLKINVX2TS U9266 ( .A(n1714), .Y(n12475) );
  INVX1TS U9267 ( .A(n10421), .Y(n10902) );
  INVX2TS U9268 ( .A(n10534), .Y(n11148) );
  CLKINVX1TS U9269 ( .A(n10440), .Y(n10931) );
  CLKINVX2TS U9270 ( .A(n5342), .Y(n12386) );
  AOI22X1TS U9271 ( .A0(n12512), .A1(n12265), .B0(n11269), .B1(n5353), .Y(
        n5688) );
  INVXLTS U9272 ( .A(n2423), .Y(n9058) );
  INVX1TS U9273 ( .A(n7651), .Y(n12361) );
  AOI22XLTS U9274 ( .A0(n12635), .A1(n12344), .B0(n11170), .B1(n12473), .Y(
        n8388) );
  CLKINVX2TS U9275 ( .A(n12325), .Y(n10695) );
  INVX2TS U9276 ( .A(n10925), .Y(n11006) );
  INVX1TS U9277 ( .A(n1675), .Y(n12563) );
  INVX2TS U9278 ( .A(n12251), .Y(n10424) );
  CLKINVX2TS U9279 ( .A(n7698), .Y(n9857) );
  CLKINVX2TS U9280 ( .A(n9933), .Y(n10938) );
  CLKINVX2TS U9281 ( .A(n10587), .Y(n11548) );
  CLKINVX2TS U9282 ( .A(n1750), .Y(n11608) );
  CLKINVX2TS U9283 ( .A(n2466), .Y(n10523) );
  CLKINVX2TS U9284 ( .A(n11628), .Y(n10609) );
  CLKINVX2TS U9285 ( .A(n3991), .Y(n10764) );
  INVX1TS U9286 ( .A(n5428), .Y(n11978) );
  INVX2TS U9287 ( .A(n7651), .Y(n12362) );
  INVX2TS U9288 ( .A(n11275), .Y(n10427) );
  INVX2TS U9289 ( .A(n12345), .Y(n11587) );
  INVX1TS U9290 ( .A(n3531), .Y(n10490) );
  INVX2TS U9291 ( .A(n12450), .Y(n10190) );
  INVX2TS U9292 ( .A(n7299), .Y(n12480) );
  INVX2TS U9293 ( .A(n7591), .Y(n12177) );
  INVX2TS U9294 ( .A(n10926), .Y(n10754) );
  CLKINVX2TS U9295 ( .A(n3486), .Y(n10164) );
  INVX1TS U9296 ( .A(n7229), .Y(n10018) );
  INVX2TS U9297 ( .A(n12028), .Y(n11680) );
  INVX1TS U9298 ( .A(n5506), .Y(n10465) );
  INVX1TS U9299 ( .A(n1675), .Y(n12564) );
  INVX1TS U9300 ( .A(n3630), .Y(n12039) );
  CLKINVX1TS U9301 ( .A(n5600), .Y(n10487) );
  CLKINVX2TS U9302 ( .A(n2466), .Y(n10524) );
  INVX2TS U9303 ( .A(n2628), .Y(n10509) );
  INVX2TS U9304 ( .A(n3544), .Y(n12443) );
  INVX1TS U9305 ( .A(n5514), .Y(n11698) );
  INVX1TS U9306 ( .A(n11145), .Y(n11109) );
  CLKINVX2TS U9307 ( .A(n10514), .Y(n11017) );
  INVX1TS U9308 ( .A(n2245), .Y(n10993) );
  INVX2TS U9309 ( .A(n11030), .Y(n11852) );
  CLKINVX2TS U9310 ( .A(n5293), .Y(n10824) );
  INVX2TS U9311 ( .A(n5298), .Y(n11689) );
  CLKINVX2TS U9312 ( .A(n11229), .Y(n10501) );
  CLKINVX2TS U9313 ( .A(n4321), .Y(n12493) );
  INVX1TS U9314 ( .A(n4501), .Y(n10812) );
  CLKINVX1TS U9315 ( .A(n3930), .Y(n12568) );
  CLKINVX2TS U9316 ( .A(n3691), .Y(n10850) );
  CLKINVX2TS U9317 ( .A(n5478), .Y(n11264) );
  CLKINVX2TS U9318 ( .A(n5761), .Y(n11373) );
  INVX1TS U9319 ( .A(n5622), .Y(n12440) );
  CLKINVX2TS U9320 ( .A(n12017), .Y(n9676) );
  CLKINVX2TS U9321 ( .A(n12074), .Y(n10503) );
  INVX1TS U9322 ( .A(n7462), .Y(n11119) );
  CLKINVX2TS U9323 ( .A(n5446), .Y(n10892) );
  CLKINVX2TS U9324 ( .A(n10734), .Y(n12322) );
  CLKINVX2TS U9325 ( .A(n12072), .Y(n10504) );
  INVX1TS U9326 ( .A(n9528), .Y(n12471) );
  INVX1TS U9327 ( .A(n3827), .Y(n12388) );
  OAI21XLTS U9328 ( .A0(n12308), .A1(n11442), .B0(n12341), .Y(n3061) );
  CLKINVX2TS U9329 ( .A(n3870), .Y(n9658) );
  CLKINVX2TS U9330 ( .A(n11057), .Y(n11948) );
  CLKINVX1TS U9331 ( .A(n1758), .Y(n10654) );
  INVX1TS U9332 ( .A(n7512), .Y(n11565) );
  INVX2TS U9333 ( .A(n3895), .Y(n9654) );
  INVX1TS U9334 ( .A(n2069), .Y(n11042) );
  INVX2TS U9335 ( .A(n1819), .Y(n12359) );
  INVX2TS U9336 ( .A(n1819), .Y(n12358) );
  NOR2X1TS U9337 ( .A(n10539), .B(n12373), .Y(n2311) );
  INVX1TS U9338 ( .A(n2291), .Y(n12086) );
  CLKINVX2TS U9339 ( .A(n2307), .Y(n10548) );
  CLKINVX2TS U9340 ( .A(n7767), .Y(n11932) );
  INVX1TS U9341 ( .A(n12139), .Y(n12176) );
  INVX2TS U9342 ( .A(n9527), .Y(n12470) );
  CLKINVX2TS U9343 ( .A(n10635), .Y(n10999) );
  INVX2TS U9344 ( .A(n11025), .Y(n11603) );
  INVX2TS U9345 ( .A(n7166), .Y(n11050) );
  CLKINVX1TS U9346 ( .A(n5798), .Y(n10985) );
  AOI22X1TS U9347 ( .A0(n11683), .A1(n12450), .B0(n10562), .B1(n11337), .Y(
        n6045) );
  CLKINVX2TS U9348 ( .A(n12145), .Y(n10208) );
  INVX1TS U9349 ( .A(n2629), .Y(n12290) );
  CLKINVX1TS U9350 ( .A(n3554), .Y(n12254) );
  INVX1TS U9351 ( .A(n7403), .Y(n11547) );
  CLKINVX2TS U9352 ( .A(n3530), .Y(n10494) );
  INVX1TS U9353 ( .A(n3762), .Y(n10816) );
  INVX1TS U9354 ( .A(n5367), .Y(n10440) );
  CLKINVX1TS U9355 ( .A(n5391), .Y(n12258) );
  CLKINVX2TS U9356 ( .A(n3649), .Y(n10867) );
  CLKINVX2TS U9357 ( .A(n1972), .Y(n10630) );
  CLKINVX1TS U9358 ( .A(n7964), .Y(n11952) );
  INVX2TS U9359 ( .A(n5484), .Y(n12265) );
  INVX1TS U9360 ( .A(n7131), .Y(n12096) );
  CLKINVX2TS U9361 ( .A(n2013), .Y(n12557) );
  INVX1TS U9362 ( .A(n7090), .Y(n11795) );
  CLKINVX2TS U9363 ( .A(n7589), .Y(n12164) );
  CLKINVX1TS U9364 ( .A(n3593), .Y(n12231) );
  INVX2TS U9365 ( .A(n3794), .Y(n11285) );
  CLKINVX2TS U9366 ( .A(n7488), .Y(n11902) );
  INVX2TS U9367 ( .A(n6012), .Y(n10555) );
  CLKINVX1TS U9368 ( .A(n7649), .Y(n12356) );
  INVX1TS U9369 ( .A(n1718), .Y(n10672) );
  INVX2TS U9370 ( .A(n3758), .Y(n12396) );
  INVX1TS U9371 ( .A(n5328), .Y(n10422) );
  CLKINVX1TS U9372 ( .A(n5352), .Y(n12235) );
  CLKINVX2TS U9373 ( .A(n5395), .Y(n12407) );
  CLKINVX2TS U9374 ( .A(n12588), .Y(n9633) );
  CLKINVX2TS U9375 ( .A(n3597), .Y(n12419) );
  CLKINVX2TS U9376 ( .A(n5356), .Y(n12391) );
  CLKINVX2TS U9377 ( .A(n7715), .Y(n9862) );
  CLKINVX1TS U9378 ( .A(n5352), .Y(n12234) );
  CLKINVX1TS U9379 ( .A(n7144), .Y(n12102) );
  CLKINVX1TS U9380 ( .A(n7313), .Y(n10286) );
  CLKINVX2TS U9381 ( .A(n3575), .Y(n10467) );
  CLKINVX2TS U9382 ( .A(n3672), .Y(n11755) );
  INVX1TS U9383 ( .A(n11298), .Y(n9910) );
  CLKINVX2TS U9384 ( .A(n7337), .Y(n11522) );
  CLKINVX1TS U9385 ( .A(n5356), .Y(n12394) );
  AOI22X1TS U9386 ( .A0(n11711), .A1(n11282), .B0(n11221), .B1(n12520), .Y(
        n5905) );
  CLKINVX2TS U9387 ( .A(n5744), .Y(n9982) );
  INVX2TS U9388 ( .A(n7086), .Y(n11783) );
  AOI22X1TS U9389 ( .A0(n11738), .A1(n11369), .B0(n11404), .B1(n12524), .Y(
        n4049) );
  INVX1TS U9390 ( .A(n1756), .Y(n10659) );
  CLKINVX2TS U9391 ( .A(n1976), .Y(n10625) );
  CLKINVX2TS U9392 ( .A(n2061), .Y(n9090) );
  INVX1TS U9393 ( .A(n2492), .Y(n10515) );
  INVX1TS U9394 ( .A(n2638), .Y(n11817) );
  INVX2TS U9395 ( .A(n12269), .Y(n9153) );
  INVX1TS U9396 ( .A(n1709), .Y(n12601) );
  INVX2TS U9397 ( .A(n1869), .Y(n12144) );
  INVX1TS U9398 ( .A(n2363), .Y(n10527) );
  CLKINVX2TS U9399 ( .A(n2141), .Y(n11835) );
  CLKINVX2TS U9400 ( .A(n2042), .Y(n10602) );
  CLKINVX2TS U9401 ( .A(n10553), .Y(n11632) );
  CLKINVX1TS U9402 ( .A(n1663), .Y(n10016) );
  CLKINVX2TS U9403 ( .A(n3672), .Y(n11756) );
  INVX1TS U9404 ( .A(n12015), .Y(n12018) );
  CLKINVX2TS U9405 ( .A(n3558), .Y(n12435) );
  CLKINVX2TS U9406 ( .A(n12584), .Y(n9636) );
  INVX2TS U9407 ( .A(n12005), .Y(n10181) );
  CLKINVX1TS U9408 ( .A(n2649), .Y(n11442) );
  CLKINVX2TS U9409 ( .A(n10688), .Y(n9817) );
  CLKINVX2TS U9410 ( .A(n3929), .Y(n12573) );
  INVX2TS U9411 ( .A(n1869), .Y(n12147) );
  CLKINVX2TS U9412 ( .A(n6094), .Y(n10567) );
  INVX1TS U9413 ( .A(n7113), .Y(n10605) );
  INVX1TS U9414 ( .A(n3820), .Y(n10801) );
  CLKINVX2TS U9415 ( .A(n7843), .Y(n11610) );
  INVX1TS U9416 ( .A(n5876), .Y(n10531) );
  CLKINVX2TS U9417 ( .A(n1887), .Y(n11888) );
  CLKINVX2TS U9418 ( .A(n3869), .Y(n11261) );
  CLKINVX2TS U9419 ( .A(n7070), .Y(n11421) );
  INVX1TS U9420 ( .A(n2480), .Y(n10962) );
  CLKINVX1TS U9421 ( .A(n7126), .Y(n12081) );
  CLKINVX1TS U9422 ( .A(n7358), .Y(n10034) );
  INVX1TS U9423 ( .A(n7648), .Y(n10062) );
  CLKINVX2TS U9424 ( .A(n5337), .Y(n12220) );
  CLKINVX2TS U9425 ( .A(n7378), .Y(n11541) );
  CLKINVX1TS U9426 ( .A(n7316), .Y(n10657) );
  CLKINVX2TS U9427 ( .A(n5337), .Y(n12218) );
  CLKINVX2TS U9428 ( .A(n5306), .Y(n12211) );
  CLKINVX2TS U9429 ( .A(n3578), .Y(n12246) );
  CLKINVX2TS U9430 ( .A(n2564), .Y(n9928) );
  INVX2TS U9431 ( .A(n7110), .Y(n12077) );
  INVX1TS U9432 ( .A(n4326), .Y(n10797) );
  INVX1TS U9433 ( .A(n1746), .Y(n12367) );
  INVX1TS U9434 ( .A(n5515), .Y(n12521) );
  INVX1TS U9435 ( .A(n3694), .Y(n12525) );
  CLKINVX2TS U9436 ( .A(n7243), .Y(n12121) );
  CLKINVX2TS U9437 ( .A(n7291), .Y(n12625) );
  CLKINVX1TS U9438 ( .A(n2019), .Y(n11058) );
  INVXLTS U9439 ( .A(n1746), .Y(n12368) );
  INVX1TS U9440 ( .A(n8192), .Y(n11641) );
  CLKINVX2TS U9441 ( .A(n4184), .Y(n10377) );
  INVX1TS U9442 ( .A(n5311), .Y(n11679) );
  CLKINVX2TS U9443 ( .A(n5663), .Y(n12004) );
  CLKINVX2TS U9444 ( .A(n5762), .Y(n11753) );
  INVX1TS U9445 ( .A(n6138), .Y(n10572) );
  INVX1TS U9446 ( .A(n1904), .Y(n10260) );
  CLKINVX2TS U9447 ( .A(n7079), .Y(n10601) );
  CLKINVX2TS U9448 ( .A(n5306), .Y(n12212) );
  CLKINVX2TS U9449 ( .A(n5369), .Y(n11216) );
  INVX1TS U9450 ( .A(n5531), .Y(n11306) );
  CLKINVX2TS U9451 ( .A(n3532), .Y(n11411) );
  CLKINVX2TS U9452 ( .A(n6013), .Y(n9743) );
  CLKINVX2TS U9453 ( .A(n5573), .Y(n10474) );
  INVX2TS U9454 ( .A(n2163), .Y(n9952) );
  CLKAND2X2TS U9455 ( .A(n7226), .B(n8600), .Y(n7126) );
  CLKINVX2TS U9456 ( .A(n2278), .Y(n9716) );
  CLKINVX2TS U9457 ( .A(n3659), .Y(n11380) );
  CLKINVX2TS U9458 ( .A(n4273), .Y(n10384) );
  AND2X2TS U9459 ( .A(n4742), .B(n4938), .Y(n3614) );
  CLKINVX2TS U9460 ( .A(n4514), .Y(n9683) );
  CLKINVX2TS U9461 ( .A(n6776), .Y(n9440) );
  CLKINVX2TS U9462 ( .A(n2121), .Y(n11839) );
  CLKINVX2TS U9463 ( .A(n5035), .Y(n9252) );
  CLKINVX2TS U9464 ( .A(n6834), .Y(n9448) );
  CLKINVX2TS U9465 ( .A(n5006), .Y(n9249) );
  CLKINVX2TS U9466 ( .A(n4246), .Y(n9653) );
  CLKINVX2TS U9467 ( .A(n2345), .Y(n9712) );
  CLKINVX2TS U9468 ( .A(n2095), .Y(n11845) );
  INVX1TS U9469 ( .A(n1727), .Y(n11137) );
  CLKINVX2TS U9470 ( .A(n6747), .Y(n9437) );
  CLKINVX2TS U9471 ( .A(n6585), .Y(n9432) );
  CLKINVX2TS U9472 ( .A(n4000), .Y(n9926) );
  CLKINVX2TS U9473 ( .A(n4806), .Y(n9236) );
  CLKINVX2TS U9474 ( .A(n2385), .Y(n9940) );
  CLKINVX2TS U9475 ( .A(n8116), .Y(n9580) );
  CLKINVX2TS U9476 ( .A(n4785), .Y(n9232) );
  CLKINVX2TS U9477 ( .A(n5821), .Y(n9986) );
  CLKINVX2TS U9478 ( .A(n8050), .Y(n9570) );
  CLKINVX2TS U9479 ( .A(n10736), .Y(n10737) );
  INVX2TS U9480 ( .A(n1769), .Y(n9119) );
  CLKINVX2TS U9481 ( .A(n11179), .Y(n11181) );
  CLKINVX2TS U9482 ( .A(n10348), .Y(n10350) );
  INVX1TS U9483 ( .A(n9442), .Y(n9443) );
  CLKINVX2TS U9484 ( .A(n1731), .Y(n9123) );
  CLKINVX2TS U9485 ( .A(n9404), .Y(n9405) );
  CLKINVX2TS U9486 ( .A(n9327), .Y(n9328) );
  CLKINVX2TS U9487 ( .A(n9567), .Y(n9568) );
  CLKINVX2TS U9488 ( .A(n9289), .Y(n9290) );
  CLKINVX2TS U9489 ( .A(n9309), .Y(n9310) );
  CLKINVX2TS U9490 ( .A(n9417), .Y(n9418) );
  CLKINVX2TS U9491 ( .A(n9517), .Y(n9518) );
  CLKINVX2TS U9492 ( .A(n9594), .Y(n9595) );
  CLKINVX2TS U9493 ( .A(n9468), .Y(n9469) );
  CLKINVX2TS U9494 ( .A(n9507), .Y(n9508) );
  CLKINVX2TS U9495 ( .A(n9331), .Y(n9332) );
  INVXLTS U9496 ( .A(n9412), .Y(n9414) );
  CLKINVX2TS U9497 ( .A(n9604), .Y(n9605) );
  INVXLTS U9498 ( .A(n9502), .Y(n9504) );
  CLKINVX2TS U9499 ( .A(n9314), .Y(n9315) );
  CLKINVX1TS U9500 ( .A(n9323), .Y(n9325) );
  CLKINVX2TS U9501 ( .A(n9408), .Y(n9409) );
  INVXLTS U9502 ( .A(n9586), .Y(n9588) );
  CLKINVX2TS U9503 ( .A(n9340), .Y(n9341) );
  CLKINVX1TS U9504 ( .A(n9497), .Y(n9499) );
  CLKINVX2TS U9505 ( .A(n9488), .Y(n9489) );
  INVXLTS U9506 ( .A(n9577), .Y(n9579) );
  CLKINVX2TS U9507 ( .A(n9399), .Y(n9400) );
  CLKINVX2TS U9508 ( .A(n9319), .Y(n9320) );
  CLKINVX2TS U9509 ( .A(n9548), .Y(n9549) );
  INVXLTS U9510 ( .A(n9493), .Y(n9495) );
  CLKINVX2TS U9511 ( .A(n9426), .Y(n9427) );
  CLKINVX2TS U9512 ( .A(n9377), .Y(n9378) );
  CLKINVX2TS U9513 ( .A(n9412), .Y(n9413) );
  CLKINVX2TS U9514 ( .A(n9599), .Y(n9600) );
  CLKINVX1TS U9515 ( .A(n9408), .Y(n9410) );
  INVXLTS U9516 ( .A(n9394), .Y(n9396) );
  CLKINVX2TS U9517 ( .A(n9394), .Y(n9395) );
  INVXLTS U9518 ( .A(n9309), .Y(n9311) );
  CLKINVX2TS U9519 ( .A(n9512), .Y(n9513) );
  CLKINVX2TS U9520 ( .A(n9304), .Y(n9305) );
  CLKINVX2TS U9521 ( .A(n9582), .Y(n9583) );
  INVXLTS U9522 ( .A(n9327), .Y(n9329) );
  CLKINVX2TS U9523 ( .A(n9389), .Y(n9390) );
  CLKINVX2TS U9524 ( .A(n9557), .Y(n9558) );
  CLKINVX2TS U9525 ( .A(n9590), .Y(n9591) );
  CLKINVX2TS U9526 ( .A(n9473), .Y(n9474) );
  CLKINVX2TS U9527 ( .A(n9577), .Y(n9578) );
  CLKINVX1TS U9528 ( .A(n9582), .Y(n9584) );
  INVXLTS U9529 ( .A(n9483), .Y(n9485) );
  INVXLTS U9530 ( .A(n9381), .Y(n9382) );
  INVXLTS U9531 ( .A(n9426), .Y(n9428) );
  INVXLTS U9532 ( .A(n9294), .Y(n9295) );
  INVX2TS U9533 ( .A(n9294), .Y(n9296) );
  INVXLTS U9534 ( .A(n9421), .Y(n9423) );
  INVXLTS U9535 ( .A(n9417), .Y(n9419) );
  CLKINVX2TS U9536 ( .A(n9385), .Y(n9386) );
  INVXLTS U9537 ( .A(n9340), .Y(n9342) );
  CLKINVX2TS U9538 ( .A(n9614), .Y(n9615) );
  CLKINVX2TS U9539 ( .A(n9299), .Y(n9300) );
  CLKINVX2TS U9540 ( .A(n9619), .Y(n9620) );
  CLKINVX2TS U9541 ( .A(n9609), .Y(n9610) );
  INVXLTS U9542 ( .A(n9331), .Y(n9333) );
  INVXLTS U9543 ( .A(n9604), .Y(n9606) );
  CLKINVX2TS U9544 ( .A(n9478), .Y(n9479) );
  INVXLTS U9545 ( .A(n9289), .Y(n9291) );
  INVXLTS U9546 ( .A(n9590), .Y(n9592) );
  INVXLTS U9547 ( .A(n9377), .Y(n9379) );
  CLKINVX1TS U9548 ( .A(n9517), .Y(n9519) );
  INVXLTS U9549 ( .A(n9548), .Y(n9550) );
  INVXLTS U9550 ( .A(n9473), .Y(n9475) );
  INVXLTS U9551 ( .A(n9299), .Y(n9301) );
  INVXLTS U9552 ( .A(n9385), .Y(n9387) );
  CLKINVX1TS U9553 ( .A(n9557), .Y(n9559) );
  CLKINVX2TS U9554 ( .A(n9421), .Y(n9422) );
  CLKINVX1TS U9555 ( .A(n9567), .Y(n9569) );
  CLKINVX2TS U9556 ( .A(n9336), .Y(n9337) );
  CLKINVX2TS U9557 ( .A(n9562), .Y(n9563) );
  CLKINVX2TS U9558 ( .A(n9572), .Y(n9573) );
  CLKINVX2TS U9559 ( .A(n9497), .Y(n9498) );
  CLKINVX2TS U9560 ( .A(n9586), .Y(n9587) );
  CLKINVX2TS U9561 ( .A(n9553), .Y(n9554) );
  INVXLTS U9562 ( .A(n9507), .Y(n9509) );
  CLKINVX2TS U9563 ( .A(n9483), .Y(n9484) );
  CLKINVX1TS U9564 ( .A(n9572), .Y(n9574) );
  INVXLTS U9565 ( .A(n9389), .Y(n9391) );
  CLKINVX1TS U9566 ( .A(n9512), .Y(n9514) );
  CLKINVX2TS U9567 ( .A(n9323), .Y(n9324) );
  CLKINVX2TS U9568 ( .A(n9502), .Y(n9503) );
  CLKINVX2TS U9569 ( .A(n9464), .Y(n9465) );
  INVXLTS U9570 ( .A(n9304), .Y(n9306) );
  INVXLTS U9571 ( .A(n9468), .Y(n9470) );
  INVXLTS U9572 ( .A(n9399), .Y(n9401) );
  CLKINVX2TS U9573 ( .A(n9493), .Y(n9494) );
  INVXLTS U9574 ( .A(w3[28]), .Y(n9604) );
  INVXLTS U9575 ( .A(w0[11]), .Y(n9309) );
  INVXLTS U9576 ( .A(w0[19]), .Y(n9323) );
  INVXLTS U9577 ( .A(w0[25]), .Y(n9331) );
  INVXLTS U9578 ( .A(w1[27]), .Y(n9421) );
  INVXLTS U9579 ( .A(w2[19]), .Y(n9497) );
  INVXLTS U9580 ( .A(w1[28]), .Y(n9426) );
  CLKINVX2TS U9581 ( .A(w1[3]), .Y(n9381) );
  INVXLTS U9582 ( .A(w1[20]), .Y(n9412) );
  CLKINVX1TS U9583 ( .A(w0[3]), .Y(n9294) );
  CLKINVX1TS U9584 ( .A(w2[12]), .Y(n9488) );
  INVXLTS U9585 ( .A(w0[9]), .Y(n9304) );
  INVXLTS U9586 ( .A(w1[9]), .Y(n9389) );
  INVXLTS U9587 ( .A(w3[4]), .Y(n9557) );
  INVXLTS U9588 ( .A(w3[25]), .Y(n9590) );
  INVXLTS U9589 ( .A(w2[4]), .Y(n9473) );
  INVXLTS U9590 ( .A(w1[11]), .Y(n9394) );
  INVXLTS U9591 ( .A(w3[17]), .Y(n9577) );
  INVXLTS U9592 ( .A(w2[27]), .Y(n9512) );
  INVXLTS U9593 ( .A(w3[19]), .Y(n9582) );
  INVXLTS U9594 ( .A(w0[20]), .Y(n9327) );
  INVX2TS U9595 ( .A(w1[4]), .Y(n9385) );
  INVX2TS U9596 ( .A(w0[4]), .Y(n9299) );
  INVX2TS U9597 ( .A(w2[28]), .Y(n9517) );
  INVXLTS U9598 ( .A(w0[1]), .Y(n9289) );
  INVX2TS U9599 ( .A(w2[25]), .Y(n9507) );
  INVXLTS U9600 ( .A(w2[20]), .Y(n9502) );
  INVXLTS U9601 ( .A(w3[20]), .Y(n9586) );
  INVXLTS U9602 ( .A(w0[28]), .Y(n9340) );
  INVX2TS U9603 ( .A(w3[12]), .Y(n9572) );
  INVXLTS U9604 ( .A(w3[1]), .Y(n9548) );
  INVX2TS U9605 ( .A(w1[1]), .Y(n9377) );
  INVXLTS U9606 ( .A(w1[12]), .Y(n9399) );
  INVXLTS U9607 ( .A(w2[3]), .Y(n9468) );
  INVXLTS U9608 ( .A(w2[17]), .Y(n9493) );
  INVXLTS U9609 ( .A(w1[25]), .Y(n9417) );
  INVX2TS U9610 ( .A(w3[11]), .Y(n9567) );
  INVX2TS U9611 ( .A(w1[19]), .Y(n9408) );
  INVX1TS U9612 ( .A(n5139), .Y(n9264) );
  INVX1TS U9613 ( .A(n5197), .Y(n9275) );
  CLKINVX2TS U9614 ( .A(n5139), .Y(n9263) );
  CLKINVX2TS U9615 ( .A(n3331), .Y(n9074) );
  INVX1TS U9616 ( .A(n2230), .Y(n9083) );
  CLKINVX2TS U9617 ( .A(n5125), .Y(n9260) );
  INVX1TS U9618 ( .A(n6965), .Y(n9219) );
  INVX1TS U9619 ( .A(n6965), .Y(n9220) );
  INVX1TS U9620 ( .A(n4024), .Y(n9126) );
  INVX1TS U9621 ( .A(n6991), .Y(n9459) );
  INVX1TS U9622 ( .A(n1361), .Y(n9777) );
  INVX1TS U9623 ( .A(n3386), .Y(n9194) );
  INVX2TS U9624 ( .A(n9772), .Y(n9773) );
  INVX1TS U9625 ( .A(n5182), .Y(n9209) );
  INVX1TS U9626 ( .A(n5140), .Y(n9206) );
  INVX1TS U9627 ( .A(n1402), .Y(n9234) );
  INVX1TS U9628 ( .A(n6980), .Y(n9127) );
  INVXLTS U9629 ( .A(n3338), .Y(n9134) );
  INVX1TS U9630 ( .A(n3338), .Y(n9133) );
  INVX1TS U9631 ( .A(n5186), .Y(n9116) );
  INVXLTS U9632 ( .A(n1594), .Y(n10024) );
  CLKINVX1TS U9633 ( .A(n7009), .Y(n9178) );
  INVX1TS U9634 ( .A(n5238), .Y(n9198) );
  CLKINVX1TS U9635 ( .A(n5238), .Y(n9199) );
  INVX1TS U9636 ( .A(n7009), .Y(n9177) );
  INVX1TS U9637 ( .A(n6924), .Y(n9155) );
  INVXLTS U9638 ( .A(n6924), .Y(n9156) );
  INVX1TS U9639 ( .A(n5124), .Y(n9142) );
  CLKINVX2TS U9640 ( .A(n1511), .Y(n9223) );
  INVX1TS U9641 ( .A(n3441), .Y(n9184) );
  INVXLTS U9642 ( .A(n5124), .Y(n9143) );
  INVX2TS U9643 ( .A(n1777), .Y(n9752) );
  CLKINVX2TS U9644 ( .A(n1370), .Y(n9250) );
  INVX1TS U9645 ( .A(n1997), .Y(n9737) );
  INVX1TS U9646 ( .A(n1615), .Y(n9769) );
  INVX1TS U9647 ( .A(n3346), .Y(n9187) );
  INVX1TS U9648 ( .A(n3390), .Y(n9101) );
  INVX1TS U9649 ( .A(n3330), .Y(n9130) );
  INVX1TS U9650 ( .A(n3390), .Y(n9100) );
  INVXLTS U9651 ( .A(n1995), .Y(n12659) );
  INVX2TS U9652 ( .A(n1626), .Y(n9139) );
  INVX2TS U9653 ( .A(n1584), .Y(n9167) );
  INVX2TS U9654 ( .A(n1312), .Y(n9273) );
  INVX1TS U9655 ( .A(n1387), .Y(n9239) );
  INVX2TS U9656 ( .A(n1570), .Y(n9173) );
  INVX2TS U9657 ( .A(n1616), .Y(n9148) );
  CLKINVX1TS U9658 ( .A(n6925), .Y(n9152) );
  INVX1TS U9659 ( .A(n6925), .Y(n9151) );
  INVX2TS U9660 ( .A(n1630), .Y(n9136) );
  INVX1TS U9661 ( .A(n1329), .Y(n9257) );
  INVX1TS U9662 ( .A(n1329), .Y(n9258) );
  CLKINVX1TS U9663 ( .A(n1595), .Y(n9164) );
  INVX1TS U9664 ( .A(n1305), .Y(n9780) );
  NOR4XLTS U9665 ( .A(n7097), .B(n7228), .C(n8036), .D(n8037), .Y(n6933) );
  CLKINVX1TS U9666 ( .A(n1623), .Y(n9146) );
  INVX1TS U9667 ( .A(n1637), .Y(n10020) );
  CLKINVX1TS U9668 ( .A(n6151), .Y(n9288) );
  AOI211XLTS U9669 ( .A0(n11512), .A1(n9087), .B0(n2974), .C0(n2178), .Y(n2972) );
  CLKINVX2TS U9670 ( .A(n6151), .Y(n9287) );
  INVX1TS U9671 ( .A(n4204), .Y(n9165) );
  INVX1TS U9672 ( .A(n6114), .Y(n9371) );
  INVX1TS U9673 ( .A(n5973), .Y(n9352) );
  INVX1TS U9674 ( .A(n6070), .Y(n9363) );
  INVX1TS U9675 ( .A(n4160), .Y(n9157) );
  CLKINVX2TS U9676 ( .A(n7359), .Y(n9826) );
  INVX2TS U9677 ( .A(n1668), .Y(n12188) );
  CLKINVX2TS U9678 ( .A(n7209), .Y(n9814) );
  CLKINVX2TS U9679 ( .A(n7067), .Y(n9798) );
  CLKINVX1TS U9680 ( .A(n7315), .Y(n10651) );
  CLKINVX2TS U9681 ( .A(n1986), .Y(n11555) );
  AOI22XLTS U9682 ( .A0(n12124), .A1(n11839), .B0(n11924), .B1(n2453), .Y(
        n2450) );
  CLKINVX2TS U9683 ( .A(n11024), .Y(n11080) );
  CLKINVX2TS U9684 ( .A(n7734), .Y(n10724) );
  INVX1TS U9685 ( .A(n2628), .Y(n10510) );
  INVX1TS U9686 ( .A(n9190), .Y(n12208) );
  INVX1TS U9687 ( .A(n7314), .Y(n10647) );
  CLKINVX2TS U9688 ( .A(n7314), .Y(n10648) );
  OAI31X1TS U9689 ( .A0(n12240), .A1(n12255), .A2(n10465), .B0(n12249), .Y(
        n5505) );
  CLKINVX2TS U9690 ( .A(n10917), .Y(n11350) );
  INVX2TS U9691 ( .A(n12266), .Y(n9703) );
  CLKINVX2TS U9692 ( .A(n10851), .Y(n11251) );
  CLKINVX2TS U9693 ( .A(n10587), .Y(n11549) );
  CLKINVX1TS U9694 ( .A(n7276), .Y(n12128) );
  INVX1TS U9695 ( .A(n2379), .Y(n9064) );
  CLKINVX2TS U9696 ( .A(n3518), .Y(n10921) );
  CLKINVX2TS U9697 ( .A(n7155), .Y(n10665) );
  INVX1TS U9698 ( .A(n10476), .Y(n10811) );
  CLKINVX2TS U9699 ( .A(n10870), .Y(n11300) );
  AOI22X1TS U9700 ( .A0(n11266), .A1(n11810), .B0(n12073), .B1(n12592), .Y(
        n4756) );
  CLKINVX2TS U9701 ( .A(n10868), .Y(n11299) );
  INVX2TS U9702 ( .A(n12274), .Y(n9707) );
  INVX1TS U9703 ( .A(n2423), .Y(n9057) );
  CLKINVX2TS U9704 ( .A(n11014), .Y(n11287) );
  INVXLTS U9705 ( .A(n2379), .Y(n9065) );
  CLKINVX2TS U9706 ( .A(n12566), .Y(n9639) );
  INVX1TS U9707 ( .A(n9989), .Y(n10829) );
  CLKINVX2TS U9708 ( .A(n2041), .Y(n10607) );
  CLKINVX2TS U9709 ( .A(n7276), .Y(n12127) );
  INVX1TS U9710 ( .A(n10494), .Y(n10839) );
  INVX1TS U9711 ( .A(n7231), .Y(n12313) );
  CLKINVX2TS U9712 ( .A(n4296), .Y(n10792) );
  INVX1TS U9713 ( .A(n3544), .Y(n12444) );
  INVX2TS U9714 ( .A(n10625), .Y(n11011) );
  CLKINVX2TS U9715 ( .A(n10003), .Y(n10004) );
  INVX2TS U9716 ( .A(n10898), .Y(n10994) );
  CLKINVX1TS U9717 ( .A(n3671), .Y(n12024) );
  INVX2TS U9718 ( .A(n5296), .Y(n9942) );
  INVX2TS U9719 ( .A(n5342), .Y(n12383) );
  INVX1TS U9720 ( .A(n7235), .Y(n12114) );
  CLKINVX2TS U9721 ( .A(n7235), .Y(n12113) );
  CLKINVX1TS U9722 ( .A(n3996), .Y(n10403) );
  CLKINVX2TS U9723 ( .A(n11323), .Y(n10444) );
  CLKINVX1TS U9724 ( .A(n3544), .Y(n12446) );
  INVX2TS U9725 ( .A(n12163), .Y(n10090) );
  CLKINVX2TS U9726 ( .A(n7122), .Y(n12462) );
  CLKINVX2TS U9727 ( .A(n11058), .Y(n11949) );
  CLKINVX2TS U9728 ( .A(n5415), .Y(n10153) );
  INVX2TS U9729 ( .A(n1811), .Y(n11918) );
  INVX2TS U9730 ( .A(n7975), .Y(n12595) );
  INVX1TS U9731 ( .A(n10093), .Y(n11134) );
  INVX2TS U9732 ( .A(n10844), .Y(n10760) );
  CLKINVX2TS U9733 ( .A(n7163), .Y(n11819) );
  CLKINVX2TS U9734 ( .A(n5782), .Y(n10979) );
  CLKINVX2TS U9735 ( .A(n10855), .Y(n10106) );
  INVX2TS U9736 ( .A(n10835), .Y(n10186) );
  CLKINVX2TS U9737 ( .A(n11032), .Y(n11071) );
  CLKINVX1TS U9738 ( .A(n3991), .Y(n10765) );
  CLKINVX2TS U9739 ( .A(n3991), .Y(n10763) );
  INVX2TS U9740 ( .A(n10933), .Y(n10124) );
  INVX2TS U9741 ( .A(n9809), .Y(n11790) );
  CLKINVX1TS U9742 ( .A(n7235), .Y(n12115) );
  CLKINVX2TS U9743 ( .A(n5953), .Y(n11020) );
  INVX2TS U9744 ( .A(n9403), .Y(n11999) );
  CLKINVX1TS U9745 ( .A(n5844), .Y(n11385) );
  CLKINVX2TS U9746 ( .A(n7396), .Y(n10293) );
  INVX1TS U9747 ( .A(n6015), .Y(n11403) );
  CLKINVX2TS U9748 ( .A(n11938), .Y(n9467) );
  INVX1TS U9749 ( .A(n11990), .Y(n10201) );
  INVX1TS U9750 ( .A(n5798), .Y(n10984) );
  INVX1TS U9751 ( .A(n5293), .Y(n10826) );
  CLKINVX1TS U9752 ( .A(n2720), .Y(n11430) );
  CLKINVX2TS U9753 ( .A(n11028), .Y(n11851) );
  INVX1TS U9754 ( .A(n1974), .Y(n11075) );
  CLKINVX2TS U9755 ( .A(n9997), .Y(n10412) );
  CLKINVX2TS U9756 ( .A(n12308), .Y(n11035) );
  CLKINVX2TS U9757 ( .A(n1938), .Y(n12348) );
  INVX1TS U9758 ( .A(n3583), .Y(n12428) );
  CLKINVX2TS U9759 ( .A(n1749), .Y(n12467) );
  CLKINVX2TS U9760 ( .A(n1702), .Y(n10675) );
  CLKINVX2TS U9761 ( .A(n1974), .Y(n11073) );
  INVX2TS U9762 ( .A(n11996), .Y(n11731) );
  INVX2TS U9763 ( .A(n2145), .Y(n11828) );
  INVX2TS U9764 ( .A(n10895), .Y(n10443) );
  CLKINVX2TS U9765 ( .A(n11280), .Y(n10472) );
  CLKINVX1TS U9766 ( .A(n2358), .Y(n12079) );
  INVX1TS U9767 ( .A(n10533), .Y(n11149) );
  CLKINVX2TS U9768 ( .A(n11033), .Y(n11072) );
  INVX1TS U9769 ( .A(n12258), .Y(n10513) );
  INVX2TS U9770 ( .A(n12026), .Y(n11682) );
  INVX2TS U9771 ( .A(n9630), .Y(n9632) );
  INVX2TS U9772 ( .A(n10816), .Y(n10774) );
  INVX1TS U9773 ( .A(n11278), .Y(n10471) );
  CLKINVX1TS U9774 ( .A(n2687), .Y(n11436) );
  INVX2TS U9775 ( .A(n3490), .Y(n11810) );
  CLKINVX2TS U9776 ( .A(n2291), .Y(n12085) );
  CLKINVX2TS U9777 ( .A(n2380), .Y(n11482) );
  INVX2TS U9778 ( .A(n11520), .Y(n10303) );
  AND2X2TS U9779 ( .A(n6702), .B(n5625), .Y(n5798) );
  CLKINVX2TS U9780 ( .A(n11508), .Y(n10291) );
  INVX1TS U9781 ( .A(n5395), .Y(n12408) );
  CLKINVX2TS U9782 ( .A(n5700), .Y(n9714) );
  OR3X1TS U9783 ( .A(sa31[5]), .B(n9374), .C(n9874), .Y(n7725) );
  CLKINVX1TS U9784 ( .A(n12269), .Y(n9154) );
  INVX2TS U9785 ( .A(n11103), .Y(n11916) );
  CLKINVX2TS U9786 ( .A(n2240), .Y(n10574) );
  CLKINVX2TS U9787 ( .A(n7131), .Y(n12095) );
  INVX2TS U9788 ( .A(n7073), .Y(n11431) );
  INVX1TS U9789 ( .A(n5511), .Y(n10469) );
  CLKINVX1TS U9790 ( .A(n5395), .Y(n12410) );
  INVX1TS U9791 ( .A(n5445), .Y(n10462) );
  AND2X2TS U9792 ( .A(n5753), .B(n6639), .Y(n5761) );
  INVX2TS U9793 ( .A(n1686), .Y(n10003) );
  CLKINVX1TS U9794 ( .A(n3597), .Y(n12422) );
  CLKINVX2TS U9795 ( .A(n3692), .Y(n12403) );
  INVX2TS U9796 ( .A(n5447), .Y(n12417) );
  INVX2TS U9797 ( .A(n11530), .Y(n10224) );
  CLKINVX2TS U9798 ( .A(n11131), .Y(n11122) );
  AND2X2TS U9799 ( .A(n6904), .B(n6639), .Y(n5953) );
  CLKINVX2TS U9800 ( .A(n3691), .Y(n10848) );
  CLKINVX1TS U9801 ( .A(n7144), .Y(n12103) );
  CLKINVX2TS U9802 ( .A(n5446), .Y(n10890) );
  INVX1TS U9803 ( .A(n5857), .Y(n10526) );
  INVX1TS U9804 ( .A(n5356), .Y(n12392) );
  CLKINVX2TS U9805 ( .A(n12219), .Y(n9359) );
  INVX1TS U9806 ( .A(n8351), .Y(n11199) );
  INVX2TS U9807 ( .A(n7285), .Y(n11092) );
  CLKINVX2TS U9808 ( .A(n1846), .Y(n10280) );
  CLKINVX2TS U9809 ( .A(n2307), .Y(n10547) );
  INVX1TS U9810 ( .A(n4057), .Y(n10399) );
  CLKINVX1TS U9811 ( .A(n12219), .Y(n9360) );
  CLKINVX2TS U9812 ( .A(n3501), .Y(n12282) );
  CLKINVX2TS U9813 ( .A(n7169), .Y(n11467) );
  CLKINVX1TS U9814 ( .A(n3558), .Y(n12438) );
  INVX1TS U9815 ( .A(n3558), .Y(n12436) );
  CLKINVX2TS U9816 ( .A(n12641), .Y(n10356) );
  CLKINVX2TS U9817 ( .A(n12242), .Y(n9367) );
  INVX1TS U9818 ( .A(n3597), .Y(n12420) );
  INVX2TS U9819 ( .A(n3758), .Y(n12398) );
  CLKINVX2TS U9820 ( .A(n7992), .Y(n10351) );
  INVX1TS U9821 ( .A(n1720), .Y(n10666) );
  CLKINVX2TS U9822 ( .A(n7182), .Y(n11842) );
  CLKINVX1TS U9823 ( .A(n5314), .Y(n10417) );
  INVX2TS U9824 ( .A(n2469), .Y(n10965) );
  INVX2TS U9825 ( .A(n12598), .Y(n9630) );
  CLKINVX2TS U9826 ( .A(n1909), .Y(n10256) );
  CLKINVX2TS U9827 ( .A(n1751), .Y(n11600) );
  INVX1TS U9828 ( .A(n3569), .Y(n10476) );
  INVX2TS U9829 ( .A(n5513), .Y(n12425) );
  CLKINVX2TS U9830 ( .A(n5725), .Y(n9718) );
  INVX2TS U9831 ( .A(n12602), .Y(n9626) );
  CLKINVX1TS U9832 ( .A(n3729), .Y(n12223) );
  CLKINVX2TS U9833 ( .A(n2240), .Y(n10575) );
  CLKINVX1TS U9834 ( .A(n1692), .Y(n11644) );
  INVX2TS U9835 ( .A(n3627), .Y(n11787) );
  OR3X1TS U9836 ( .A(n10080), .B(sa22[6]), .C(n9252), .Y(n3597) );
  CLKINVX1TS U9837 ( .A(n3593), .Y(n12229) );
  INVX1TS U9838 ( .A(n2034), .Y(n10232) );
  CLKINVX1TS U9839 ( .A(n3752), .Y(n10828) );
  CLKINVX1TS U9840 ( .A(n7592), .Y(n12345) );
  CLKINVX2TS U9841 ( .A(n2065), .Y(n12317) );
  CLKINVX1TS U9842 ( .A(n7592), .Y(n12344) );
  INVX1TS U9843 ( .A(n5423), .Y(n11670) );
  CLKINVX2TS U9844 ( .A(n11490), .Y(n10544) );
  INVX1TS U9845 ( .A(n2196), .Y(n11005) );
  CLKINVX2TS U9846 ( .A(n5744), .Y(n9981) );
  INVX1TS U9847 ( .A(n5451), .Y(n10897) );
  CLKINVX2TS U9848 ( .A(n12002), .Y(n9668) );
  INVX1TS U9849 ( .A(n5301), .Y(n10834) );
  INVX1TS U9850 ( .A(n5294), .Y(n12196) );
  INVX1TS U9851 ( .A(n5309), .Y(n11207) );
  CLKINVX2TS U9852 ( .A(n2042), .Y(n10603) );
  CLKINVX2TS U9853 ( .A(n4081), .Y(n11996) );
  INVX2TS U9854 ( .A(n5290), .Y(n11696) );
  INVX1TS U9855 ( .A(n2952), .Y(n11422) );
  INVX2TS U9856 ( .A(n7155), .Y(n10612) );
  AND2X2TS U9857 ( .A(n5033), .B(n5040), .Y(n3758) );
  CLKINVX2TS U9858 ( .A(n7986), .Y(n10094) );
  INVX1TS U9859 ( .A(n1882), .Y(n10264) );
  CLKINVX2TS U9860 ( .A(n5724), .Y(n11366) );
  CLKINVX1TS U9861 ( .A(n3593), .Y(n12230) );
  CLKINVX1TS U9862 ( .A(n2158), .Y(n11029) );
  INVX1TS U9863 ( .A(n4076), .Y(n10394) );
  CLKINVX2TS U9864 ( .A(n7208), .Y(n9810) );
  CLKINVX1TS U9865 ( .A(n12649), .Y(n12652) );
  CLKINVX2TS U9866 ( .A(n5825), .Y(n12028) );
  CLKINVX2TS U9867 ( .A(n12202), .Y(n10775) );
  INVX2TS U9868 ( .A(n5584), .Y(n10940) );
  CLKINVX2TS U9869 ( .A(n6337), .Y(n9403) );
  INVX1TS U9870 ( .A(n5517), .Y(n10924) );
  INVX1TS U9871 ( .A(n5423), .Y(n11669) );
  CLKINVX1TS U9872 ( .A(n5391), .Y(n12257) );
  CLKINVX2TS U9873 ( .A(n5663), .Y(n12006) );
  AND2X2TS U9874 ( .A(n4975), .B(n4982), .Y(n3692) );
  INVX1TS U9875 ( .A(n5441), .Y(n10884) );
  CLKINVX2TS U9876 ( .A(n11494), .Y(n10569) );
  CLKINVX1TS U9877 ( .A(n5954), .Y(n10225) );
  INVX2TS U9878 ( .A(n5425), .Y(n11676) );
  INVX1TS U9879 ( .A(n7545), .Y(n10325) );
  INVX1TS U9880 ( .A(n5881), .Y(n12041) );
  INVX1TS U9881 ( .A(n5932), .Y(n10542) );
  CLKINVX2TS U9882 ( .A(n7244), .Y(n10628) );
  INVX2TS U9883 ( .A(n7488), .Y(n11904) );
  CLKINVX1TS U9884 ( .A(n12202), .Y(n10777) );
  CLKINVX1TS U9885 ( .A(n8477), .Y(n9874) );
  INVX1TS U9886 ( .A(n3821), .Y(n11274) );
  INVX1TS U9887 ( .A(n3503), .Y(n10932) );
  INVX1TS U9888 ( .A(n7140), .Y(n11451) );
  CLKINVX2TS U9889 ( .A(n12036), .Y(n9770) );
  INVX1TS U9890 ( .A(n3511), .Y(n11417) );
  INVX1TS U9891 ( .A(n5507), .Y(n10912) );
  INVX1TS U9892 ( .A(n5507), .Y(n10914) );
  INVX1TS U9893 ( .A(n12649), .Y(n12653) );
  OR3X1TS U9894 ( .A(n10052), .B(sa11[6]), .C(n9244), .Y(n3558) );
  CLKINVX2TS U9895 ( .A(n7109), .Y(n12306) );
  AND2X2TS U9896 ( .A(n6774), .B(n6781), .Y(n5447) );
  OR3X1TS U9897 ( .A(n10100), .B(sa23[6]), .C(n9448), .Y(n5395) );
  CLKINVX2TS U9898 ( .A(n8477), .Y(n9873) );
  CLKINVX2TS U9899 ( .A(n7243), .Y(n12119) );
  CLKINVX2TS U9900 ( .A(n5306), .Y(n12210) );
  CLKINVX1TS U9901 ( .A(n2952), .Y(n11424) );
  INVX1TS U9902 ( .A(n3686), .Y(n10854) );
  CLKINVX1TS U9903 ( .A(n3686), .Y(n10856) );
  AND2X2TS U9904 ( .A(n6832), .B(n6839), .Y(n5513) );
  CLKINVX1TS U9905 ( .A(n2296), .Y(n10557) );
  CLKINVX2TS U9906 ( .A(n2484), .Y(n11460) );
  CLKINVX1TS U9907 ( .A(n11116), .Y(n11573) );
  CLKINVX2TS U9908 ( .A(n2065), .Y(n12318) );
  CLKINVX1TS U9909 ( .A(n2158), .Y(n11030) );
  INVX1TS U9910 ( .A(n1945), .Y(n10240) );
  OR3X1TS U9911 ( .A(n10072), .B(sa12[6]), .C(n9440), .Y(n5356) );
  INVX1TS U9912 ( .A(n5441), .Y(n10886) );
  CLKINVX1TS U9913 ( .A(n5352), .Y(n12233) );
  CLKINVX2TS U9914 ( .A(n7120), .Y(n10006) );
  AND2X2TS U9915 ( .A(n4985), .B(n4975), .Y(n3869) );
  INVX1TS U9916 ( .A(n7731), .Y(n9849) );
  AND2X2TS U9917 ( .A(n3313), .B(n3321), .Y(n2484) );
  CLKINVX2TS U9918 ( .A(n7586), .Y(n12156) );
  AND2X2TS U9919 ( .A(n4876), .B(n4334), .Y(n3666) );
  AND2X2TS U9920 ( .A(n9205), .B(n4517), .Y(n3929) );
  CLKINVX2TS U9921 ( .A(n7658), .Y(n10706) );
  INVX1TS U9922 ( .A(n2188), .Y(n11518) );
  INVX1TS U9923 ( .A(n7731), .Y(n9850) );
  OR3X1TS U9924 ( .A(n10367), .B(n9225), .C(sa33[2]), .Y(n3511) );
  AND2X2TS U9925 ( .A(n8470), .B(n10078), .Y(n7337) );
  AND2X2TS U9926 ( .A(n4976), .B(n9183), .Y(n3696) );
  OR3X1TS U9927 ( .A(n9884), .B(n10742), .C(n9653), .Y(n3503) );
  INVX1TS U9928 ( .A(n2217), .Y(n9721) );
  INVX2TS U9929 ( .A(n3924), .Y(n12015) );
  CLKINVX1TS U9930 ( .A(n7658), .Y(n10707) );
  INVX1TS U9931 ( .A(n3687), .Y(n11369) );
  INVX1TS U9932 ( .A(n2198), .Y(n11823) );
  AND2X2TS U9933 ( .A(n2668), .B(n3316), .Y(n2065) );
  OR3X1TS U9934 ( .A(n9537), .B(n9444), .C(sa23[2]), .Y(n5391) );
  CLKINVX1TS U9935 ( .A(n7162), .Y(n11463) );
  CLKINVX1TS U9936 ( .A(n2189), .Y(n11514) );
  CLKINVX1TS U9937 ( .A(n3687), .Y(n11370) );
  AND2X2TS U9938 ( .A(n5034), .B(n9186), .Y(n3762) );
  INVX1TS U9939 ( .A(n3492), .Y(n12073) );
  OR3X1TS U9940 ( .A(n10753), .B(sa33[5]), .C(n9695), .Y(n3625) );
  CLKINVX1TS U9941 ( .A(n5442), .Y(n11235) );
  AND2X2TS U9942 ( .A(n6542), .B(n6737), .Y(n5412) );
  INVX2TS U9943 ( .A(n3512), .Y(n11797) );
  INVX1TS U9944 ( .A(n5311), .Y(n11677) );
  CLKINVX2TS U9945 ( .A(n5764), .Y(n12020) );
  INVX1TS U9946 ( .A(n5345), .Y(n12581) );
  INVX1TS U9947 ( .A(n5633), .Y(n10958) );
  AND2X2TS U9948 ( .A(n6784), .B(n6774), .Y(n5699) );
  OR3X1TS U9949 ( .A(sa12[3]), .B(n9836), .C(n9322), .Y(n5441) );
  INVX1TS U9950 ( .A(n3586), .Y(n12578) );
  INVX1TS U9951 ( .A(n4228), .Y(n10373) );
  CLKINVX1TS U9952 ( .A(n4256), .Y(n10374) );
  CLKINVX2TS U9953 ( .A(n5959), .Y(n10230) );
  INVX1TS U9954 ( .A(n5442), .Y(n11234) );
  CLKINVX2TS U9955 ( .A(n5574), .Y(n9711) );
  AND2X2TS U9956 ( .A(n6775), .B(n9380), .Y(n5451) );
  AND2X2TS U9957 ( .A(n6905), .B(n6674), .Y(n5663) );
  OR3X1TS U9958 ( .A(sa22[3]), .B(sa22[0]), .C(n9141), .Y(n3752) );
  INVX2TS U9959 ( .A(n5574), .Y(n9710) );
  INVX2TS U9960 ( .A(n2432), .Y(n11465) );
  CLKINVX2TS U9961 ( .A(n5760), .Y(n10518) );
  OR3X1TS U9962 ( .A(n9882), .B(n7630), .C(n10068), .Y(n7592) );
  CLKINVX1TS U9963 ( .A(n2189), .Y(n11512) );
  INVX2TS U9964 ( .A(n2198), .Y(n11821) );
  INVX1TS U9965 ( .A(n3547), .Y(n12585) );
  AND2X2TS U9966 ( .A(n8425), .B(n8479), .Y(n7843) );
  INVX1TS U9967 ( .A(n7072), .Y(n11425) );
  AND2X2TS U9968 ( .A(n6724), .B(n6737), .Y(n5306) );
  INVX1TS U9969 ( .A(n3513), .Y(n11791) );
  INVX1TS U9970 ( .A(n3665), .Y(n11376) );
  OR3X1TS U9971 ( .A(n10360), .B(n10364), .C(n3026), .Y(n2649) );
  AND2X2TS U9972 ( .A(n4876), .B(n9256), .Y(n3672) );
  INVX1TS U9973 ( .A(n5345), .Y(n12583) );
  AND2X2TS U9974 ( .A(n5106), .B(n9256), .Y(n3640) );
  INVX1TS U9975 ( .A(n3665), .Y(n11375) );
  AND2X2TS U9976 ( .A(n4517), .B(n5092), .Y(n3915) );
  INVX1TS U9977 ( .A(n3665), .Y(n11374) );
  AND2X2TS U9978 ( .A(n5043), .B(n5033), .Y(n3894) );
  INVX1TS U9979 ( .A(n4481), .Y(n12619) );
  INVX1TS U9980 ( .A(n1943), .Y(n10636) );
  INVX1TS U9981 ( .A(n3586), .Y(n12579) );
  OR3X1TS U9982 ( .A(n9434), .B(n9437), .C(n11186), .Y(n5352) );
  INVX1TS U9983 ( .A(n3838), .Y(n10794) );
  AND2X2TS U9984 ( .A(n6842), .B(n6855), .Y(n5932) );
  INVX1TS U9985 ( .A(n7280), .Y(n12637) );
  INVX1TS U9986 ( .A(n5384), .Y(n12589) );
  CLKINVX2TS U9987 ( .A(n7124), .Y(n11802) );
  INVX1TS U9988 ( .A(n7162), .Y(n11462) );
  INVX1TS U9989 ( .A(n3586), .Y(n12580) );
  CLKINVX2TS U9990 ( .A(n2164), .Y(n11532) );
  OR3X1TS U9991 ( .A(n9120), .B(n2113), .C(n9717), .Y(n2296) );
  INVX1TS U9992 ( .A(n7560), .Y(n10682) );
  AND2X2TS U9993 ( .A(n6842), .B(n6832), .Y(n5724) );
  INVX2TS U9994 ( .A(n3539), .Y(n12267) );
  AND2X2TS U9995 ( .A(n4985), .B(n4998), .Y(n4076) );
  OR3X1TS U9996 ( .A(n9124), .B(n2087), .C(n9713), .Y(n2363) );
  OR3X1TS U9997 ( .A(n9530), .B(n10096), .C(n9042), .Y(n2158) );
  INVX1TS U9998 ( .A(n8578), .Y(n9524) );
  CLKINVX2TS U9999 ( .A(n7366), .Y(n11874) );
  AND2X2TS U10000 ( .A(n2914), .B(n2410), .Y(n1838) );
  INVX2TS U10001 ( .A(n5376), .Y(n12240) );
  INVX1TS U10002 ( .A(n8578), .Y(n9523) );
  OR3X1TS U10003 ( .A(n9450), .B(n9249), .C(n11191), .Y(n3593) );
  CLKINVX2TS U10004 ( .A(n7326), .Y(n11103) );
  OR3X1TS U10005 ( .A(n10715), .B(n9820), .C(n9786), .Y(n5423) );
  OR3X1TS U10006 ( .A(sa11[3]), .B(n9828), .C(n9129), .Y(n3686) );
  OR3X1TS U10007 ( .A(n10349), .B(n3139), .C(n9056), .Y(n2952) );
  INVX2TS U10008 ( .A(n7135), .Y(n11808) );
  CLKINVX1TS U10009 ( .A(n5615), .Y(n10953) );
  CLKINVX2TS U10010 ( .A(n7548), .Y(n11129) );
  INVX1TS U10011 ( .A(n8679), .Y(n9505) );
  INVX2TS U10012 ( .A(n7134), .Y(n10265) );
  CLKINVX2TS U10013 ( .A(n7397), .Y(n12330) );
  INVX1TS U10014 ( .A(n5508), .Y(n11282) );
  INVX2TS U10015 ( .A(n2611), .Y(n10167) );
  INVX2TS U10016 ( .A(n7080), .Y(n9801) );
  AND2X2TS U10017 ( .A(n6833), .B(n9384), .Y(n5517) );
  CLKINVX1TS U10018 ( .A(n7059), .Y(n11027) );
  CLKINVX2TS U10019 ( .A(n7366), .Y(n11872) );
  CLKINVX1TS U10020 ( .A(n6024), .Y(n10558) );
  OR3X1TS U10021 ( .A(sa23[3]), .B(n9880), .C(n9339), .Y(n5507) );
  INVX1TS U10022 ( .A(n4807), .Y(n10138) );
  INVX1TS U10023 ( .A(n1981), .Y(n12623) );
  CLKINVX2TS U10024 ( .A(n7378), .Y(n11540) );
  CLKINVX2TS U10025 ( .A(n7124), .Y(n11801) );
  INVX2TS U10026 ( .A(n7135), .Y(n11807) );
  INVX1TS U10027 ( .A(n7318), .Y(n11511) );
  AND2X2TS U10028 ( .A(n2838), .B(n2454), .Y(n1901) );
  OR3X1TS U10029 ( .A(n10326), .B(n6534), .C(n9816), .Y(n5309) );
  INVX1TS U10030 ( .A(n7902), .Y(n10735) );
  OR3X1TS U10031 ( .A(n9808), .B(n10710), .C(n9743), .Y(n5301) );
  CLKINVX2TS U10032 ( .A(n7700), .Y(n10719) );
  OR3X1TS U10033 ( .A(n9350), .B(n9241), .C(sa11[2]), .Y(n3554) );
  INVX1TS U10034 ( .A(n7059), .Y(n11026) );
  CLKINVX1TS U10035 ( .A(n2236), .Y(n10580) );
  INVX1TS U10036 ( .A(n1987), .Y(n12099) );
  INVX1TS U10037 ( .A(n5895), .Y(n12049) );
  OR3X1TS U10038 ( .A(n11169), .B(n9211), .C(n9214), .Y(n3687) );
  INVX2TS U10039 ( .A(n5839), .Y(n12036) );
  INVX1TS U10040 ( .A(n5839), .Y(n12034) );
  OR3X1TS U10041 ( .A(n9876), .B(n9872), .C(n8598), .Y(n7113) );
  INVX2TS U10042 ( .A(n1908), .Y(n10641) );
  OR3X1TS U10043 ( .A(n11191), .B(n9218), .C(n9221), .Y(n3753) );
  OR3X1TS U10044 ( .A(n9860), .B(n10737), .C(n9570), .Y(n7234) );
  OR3X1TS U10045 ( .A(n10715), .B(n9820), .C(n9432), .Y(n5615) );
  AND2X2TS U10046 ( .A(n8600), .B(n8601), .Y(n7366) );
  INVX1TS U10047 ( .A(n7230), .Y(n12640) );
  OR3X1TS U10048 ( .A(n11169), .B(n9211), .C(n4993), .Y(n3547) );
  INVX1TS U10049 ( .A(n5330), .Y(n11205) );
  OR3X1TS U10050 ( .A(n11202), .B(n9420), .C(n6850), .Y(n5384) );
  AND2X2TS U10051 ( .A(n8579), .B(n8590), .Y(n7560) );
  OR3X1TS U10052 ( .A(n10044), .B(sa30[1]), .C(n9986), .Y(n5311) );
  AND2X2TS U10053 ( .A(n6901), .B(n6319), .Y(n5764) );
  INVX1TS U10054 ( .A(n8665), .Y(n10001) );
  INVX2TS U10055 ( .A(n9694), .Y(n9695) );
  AND2X2TS U10056 ( .A(n8668), .B(n8676), .Y(n7079) );
  INVX1TS U10057 ( .A(n2095), .Y(n11846) );
  INVX1TS U10058 ( .A(n3673), .Y(n12532) );
  OR3X1TS U10059 ( .A(n11185), .B(n9411), .C(n9415), .Y(n5442) );
  CLKINVX2TS U10060 ( .A(n2898), .Y(n9053) );
  INVX1TS U10061 ( .A(n6288), .Y(n11760) );
  CLKINVX1TS U10062 ( .A(n2864), .Y(n9076) );
  INVX1TS U10063 ( .A(n7158), .Y(n11814) );
  OR3X1TS U10064 ( .A(sa10[5]), .B(sa10[7]), .C(n3250), .Y(n2277) );
  OR3X1TS U10065 ( .A(n11202), .B(n9420), .C(n9424), .Y(n5508) );
  CLKINVX2TS U10066 ( .A(n2822), .Y(n9050) );
  INVX1TS U10067 ( .A(n2540), .Y(n11453) );
  INVX1TS U10068 ( .A(n6637), .Y(n9738) );
  INVX1TS U10069 ( .A(n2095), .Y(n11847) );
  AND2X2TS U10070 ( .A(n8667), .B(n8668), .Y(n7378) );
  AND2X2TS U10071 ( .A(n6910), .B(n6914), .Y(n5599) );
  OR3X1TS U10072 ( .A(sa30[0]), .B(n10709), .C(n9790), .Y(n6024) );
  INVX1TS U10073 ( .A(n4095), .Y(n11986) );
  CLKINVX2TS U10074 ( .A(n5673), .Y(n11735) );
  CLKINVX2TS U10075 ( .A(n2864), .Y(n9075) );
  OR3X1TS U10076 ( .A(sa21[5]), .B(sa21[7]), .C(n3190), .Y(n2344) );
  CLKINVX2TS U10077 ( .A(n8641), .Y(n9618) );
  OR3X1TS U10078 ( .A(n11186), .B(n9411), .C(n6792), .Y(n5345) );
  INVX1TS U10079 ( .A(n8640), .Y(n9613) );
  OR3X1TS U10080 ( .A(n3139), .B(n9696), .C(n10350), .Y(n2188) );
  CLKINVX2TS U10081 ( .A(n2121), .Y(n11840) );
  AND2X2TS U10082 ( .A(n6719), .B(n6720), .Y(n5633) );
  INVXLTS U10083 ( .A(n2540), .Y(n11454) );
  OR3X1TS U10084 ( .A(sa20[7]), .B(sa20[5]), .C(n8664), .Y(n7059) );
  AND2X2TS U10085 ( .A(n7154), .B(n8676), .Y(n7070) );
  CLKINVX2TS U10086 ( .A(n3673), .Y(n12533) );
  INVX2TS U10087 ( .A(n3776), .Y(n11297) );
  INVXLTS U10088 ( .A(n2303), .Y(n10552) );
  OR3X1TS U10089 ( .A(n9832), .B(sa02[5]), .C(n8523), .Y(n7280) );
  AND4X1TS U10090 ( .A(n8467), .B(n9585), .C(n9603), .D(n9373), .Y(n7658) );
  OR3X1TS U10091 ( .A(n10747), .B(sa33[1]), .C(n9926), .Y(n3513) );
  INVX1TS U10092 ( .A(n4273), .Y(n10386) );
  INVX1TS U10093 ( .A(n7454), .Y(n9476) );
  CLKINVX1TS U10094 ( .A(n2303), .Y(n10553) );
  AND2X2TS U10095 ( .A(n3130), .B(n2194), .Y(n1674) );
  OR3X1TS U10096 ( .A(n9193), .B(n4516), .C(sa00[2]), .Y(n3665) );
  INVX1TS U10097 ( .A(n8665), .Y(n10002) );
  OR3X1TS U10098 ( .A(n9193), .B(n5115), .C(n9788), .Y(n4481) );
  OR3X1TS U10099 ( .A(sa33[0]), .B(n10743), .C(n9699), .Y(n4256) );
  CLKINVX1TS U10100 ( .A(n2236), .Y(n10579) );
  INVX1TS U10101 ( .A(n7454), .Y(n9477) );
  INVX2TS U10102 ( .A(n3710), .Y(n11345) );
  INVX1TS U10103 ( .A(n3571), .Y(n11400) );
  AND2X2TS U10104 ( .A(n8648), .B(n9622), .Y(n7081) );
  OR3X1TS U10105 ( .A(n10752), .B(n9896), .C(n9232), .Y(n3820) );
  CLKINVX2TS U10106 ( .A(n7967), .Y(n9878) );
  CLKINVX1TS U10107 ( .A(n2940), .Y(n9069) );
  AND2X2TS U10108 ( .A(n7226), .B(n8611), .Y(n7124) );
  AND2X2TS U10109 ( .A(n8545), .B(n8535), .Y(n7586) );
  AND2X2TS U10110 ( .A(n4920), .B(n4921), .Y(n3838) );
  INVX1TS U10111 ( .A(n8599), .Y(n10262) );
  INVX1TS U10112 ( .A(n6637), .Y(n9739) );
  AND2X2TS U10113 ( .A(n8601), .B(n8611), .Y(n7133) );
  CLKINVX1TS U10114 ( .A(n4273), .Y(n10385) );
  INVX2TS U10115 ( .A(n9785), .Y(n9786) );
  CLKINVX2TS U10116 ( .A(n2940), .Y(n9068) );
  INVX1TS U10117 ( .A(n3499), .Y(n12547) );
  OR3X1TS U10118 ( .A(sa20[0]), .B(n10704), .C(n9580), .Y(n7162) );
  OR3X1TS U10119 ( .A(n11190), .B(n9218), .C(n5051), .Y(n3586) );
  INVX1TS U10120 ( .A(n8004), .Y(n11956) );
  AND2X2TS U10121 ( .A(n6911), .B(n6910), .Y(n5760) );
  INVX1TS U10122 ( .A(n7230), .Y(n12639) );
  OR3X1TS U10123 ( .A(n9525), .B(n3325), .C(n10092), .Y(n1981) );
  CLKINVX2TS U10124 ( .A(n12745), .Y(n12695) );
  AND2X2TS U10125 ( .A(n8520), .B(n9894), .Y(n8220) );
  OR3X1TS U10126 ( .A(n9461), .B(n2599), .C(n3125), .Y(n2189) );
  OR3X1TS U10127 ( .A(n9443), .B(n9439), .C(n6785), .Y(n5491) );
  CLKINVX2TS U10128 ( .A(n6420), .Y(n9416) );
  OR3X1TS U10129 ( .A(sa13[7]), .B(sa13[5]), .C(n8591), .Y(n7230) );
  CLKINVX2TS U10130 ( .A(n6420), .Y(n9415) );
  AND2X2TS U10131 ( .A(n6793), .B(n6425), .Y(n5330) );
  OR3X1TS U10132 ( .A(n10721), .B(sa01[5]), .C(n6872), .Y(n6288) );
  OR3X1TS U10133 ( .A(n11162), .B(n10309), .C(n5110), .Y(n3635) );
  OR3X1TS U10134 ( .A(sa31[5]), .B(sa31[7]), .C(n8466), .Y(n8004) );
  AND2X2TS U10135 ( .A(n6901), .B(n6910), .Y(n5573) );
  CLKINVX2TS U10136 ( .A(n2029), .Y(n9733) );
  AND2X2TS U10137 ( .A(n6910), .B(n6891), .Y(n5673) );
  OR3X1TS U10138 ( .A(n10753), .B(n9896), .C(n4929), .Y(n4273) );
  INVX2TS U10139 ( .A(n7106), .Y(n10258) );
  OR3X1TS U10140 ( .A(n10088), .B(n9848), .C(n3128), .Y(n2540) );
  AND2X2TS U10141 ( .A(n4975), .B(n4976), .Y(n3710) );
  CLKINVX2TS U10142 ( .A(n6492), .Y(n9425) );
  OR3X1TS U10143 ( .A(sa23[7]), .B(n9541), .C(n6843), .Y(n5557) );
  CLKINVX2TS U10144 ( .A(n6492), .Y(n9424) );
  AND2X2TS U10145 ( .A(n6851), .B(n6497), .Y(n5369) );
  OR3X1TS U10146 ( .A(n10032), .B(n10323), .C(n3246), .Y(n2121) );
  INVX2TS U10147 ( .A(n6564), .Y(n9785) );
  OR3X1TS U10148 ( .A(sa21[5]), .B(n10331), .C(n3184), .Y(n2303) );
  AND2X2TS U10149 ( .A(n6832), .B(n6833), .Y(n5531) );
  AND2X2TS U10150 ( .A(n8535), .B(n8520), .Y(n7611) );
  AND2X2TS U10151 ( .A(n5052), .B(n4697), .Y(n3571) );
  AND2X2TS U10152 ( .A(n4994), .B(n4625), .Y(n3532) );
  CLKINVX2TS U10153 ( .A(n4692), .Y(n9222) );
  OR3X1TS U10154 ( .A(sa22[7]), .B(n9454), .C(n5044), .Y(n3802) );
  CLKINVX2TS U10155 ( .A(n4692), .Y(n9221) );
  CLKINVX2TS U10156 ( .A(n4620), .Y(n9214) );
  OR3X1TS U10157 ( .A(sa11[7]), .B(n9355), .C(n4986), .Y(n3736) );
  CLKINVX2TS U10158 ( .A(n4620), .Y(n9215) );
  AND2X2TS U10159 ( .A(n5033), .B(n5034), .Y(n3776) );
  OR3X1TS U10160 ( .A(n9530), .B(n10096), .C(n3303), .Y(n2144) );
  INVX2TS U10161 ( .A(n4764), .Y(n9694) );
  OR3X1TS U10162 ( .A(n10032), .B(sa10[7]), .C(n3244), .Y(n2236) );
  AND2X2TS U10163 ( .A(n6774), .B(n6775), .Y(n5465) );
  OR3X1TS U10164 ( .A(n9804), .B(n9800), .C(n8657), .Y(n7158) );
  OR3X1TS U10165 ( .A(n10064), .B(n10331), .C(n3186), .Y(n2095) );
  INVX2TS U10166 ( .A(n9900), .Y(n10362) );
  INVX2TS U10167 ( .A(n11648), .Y(n11667) );
  INVX2TS U10168 ( .A(n11655), .Y(n11964) );
  INVX2TS U10169 ( .A(n11655), .Y(n11658) );
  INVX2TS U10170 ( .A(n11959), .Y(n11961) );
  INVX2TS U10171 ( .A(n11966), .Y(n11968) );
  INVX2TS U10172 ( .A(n11662), .Y(n11963) );
  INVX2TS U10173 ( .A(n11966), .Y(n11969) );
  INVX2TS U10174 ( .A(n11959), .Y(n11960) );
  INVX2TS U10175 ( .A(n11959), .Y(n11965) );
  INVX2TS U10176 ( .A(n11959), .Y(n11962) );
  INVX2TS U10177 ( .A(n11966), .Y(n11967) );
  INVX2TS U10178 ( .A(n11662), .Y(n11661) );
  INVX2TS U10179 ( .A(n11648), .Y(n11651) );
  INVX2TS U10180 ( .A(n9900), .Y(n12608) );
  CLKINVX2TS U10181 ( .A(n11173), .Y(n11175) );
  INVX2TS U10182 ( .A(n9859), .Y(n9860) );
  CLKINVX2TS U10183 ( .A(n10730), .Y(n10732) );
  CLKINVX2TS U10184 ( .A(n7656), .Y(n9854) );
  INVX1TS U10185 ( .A(n10698), .Y(n10700) );
  INVX1TS U10186 ( .A(n10725), .Y(n10727) );
  INVX2TS U10187 ( .A(n12612), .Y(n11655) );
  INVX2TS U10188 ( .A(n12612), .Y(n11959) );
  INVX2TS U10189 ( .A(n12611), .Y(n11966) );
  INVX2TS U10190 ( .A(n12611), .Y(n11662) );
  INVX2TS U10191 ( .A(n12612), .Y(n11648) );
  INVX2TS U10192 ( .A(n12606), .Y(n9900) );
  INVX2TS U10193 ( .A(sa02[2]), .Y(n10067) );
  INVX2TS U10194 ( .A(sa22[3]), .Y(n9446) );
  INVX2TS U10195 ( .A(sa31[3]), .Y(n9369) );
  INVX2TS U10196 ( .A(sa12[0]), .Y(n9835) );
  INVX2TS U10197 ( .A(sa33[2]), .Y(n9891) );
  INVX2TS U10198 ( .A(sa02[7]), .Y(n9831) );
  INVX2TS U10199 ( .A(sa33[4]), .Y(n10367) );
  INVX2TS U10200 ( .A(sa00[7]), .Y(n10317) );
  INVX2TS U10201 ( .A(sa23[4]), .Y(n9537) );
  INVX2TS U10202 ( .A(sa23[0]), .Y(n9879) );
  INVX2TS U10203 ( .A(sa22[5]), .Y(n9453) );
  INVX2TS U10204 ( .A(sa12[3]), .Y(n9430) );
  INVX2TS U10205 ( .A(sa11[0]), .Y(n9827) );
  INVX2TS U10206 ( .A(sa11[3]), .Y(n9347) );
  INVX2TS U10207 ( .A(sa30[4]), .Y(n10326) );
  INVX2TS U10208 ( .A(sa30[2]), .Y(n9815) );
  INVX2TS U10209 ( .A(sa11[5]), .Y(n9354) );
  INVX2TS U10210 ( .A(sa33[0]), .Y(n9883) );
  INVX2TS U10211 ( .A(sa22[7]), .Y(n9457) );
  INVX2TS U10212 ( .A(sa11[7]), .Y(n9357) );
  INVX2TS U10213 ( .A(sa21[1]), .Y(n9361) );
  INVX2TS U10214 ( .A(sa01[3]), .Y(n10047) );
  INVX2TS U10215 ( .A(sa33[1]), .Y(n9887) );
  INVX2TS U10216 ( .A(sa33[5]), .Y(n9895) );
  INVX2TS U10217 ( .A(sa00[3]), .Y(n10307) );
  INVX2TS U10218 ( .A(sa11[6]), .Y(n10055) );
  INVX2TS U10219 ( .A(sa31[4]), .Y(n10334) );
  INVX2TS U10220 ( .A(sa23[1]), .Y(n10099) );
  INVX2TS U10221 ( .A(sa11[1]), .Y(n10051) );
  INVX2TS U10222 ( .A(sa11[4]), .Y(n9350) );
  INVX2TS U10223 ( .A(sa21[5]), .Y(n10063) );
  INVX2TS U10224 ( .A(sa12[5]), .Y(n9438) );
  INVX2TS U10225 ( .A(sa31[6]), .Y(n10339) );
  INVX2TS U10226 ( .A(sa00[6]), .Y(n10312) );
  INVX2TS U10227 ( .A(sa30[1]), .Y(n9811) );
  INVX2TS U10228 ( .A(sa10[1]), .Y(n9281) );
  INVX2TS U10229 ( .A(sa23[3]), .Y(n9533) );
  INVX2TS U10230 ( .A(sa10[5]), .Y(n10031) );
  INVX2TS U10231 ( .A(sa12[4]), .Y(n9434) );
  INVX2TS U10232 ( .A(sa10[7]), .Y(n10322) );
  INVX2TS U10233 ( .A(sa23[6]), .Y(n10103) );
  INVX2TS U10234 ( .A(sa31[1]), .Y(n9365) );
  INVX2TS U10235 ( .A(sa30[6]), .Y(n10043) );
  INVX2TS U10236 ( .A(sa01[1]), .Y(n9823) );
  INVX2TS U10237 ( .A(sa10[3]), .Y(n10027) );
  INVX2TS U10238 ( .A(sa12[1]), .Y(n10071) );
  INVX2TS U10239 ( .A(sa22[6]), .Y(n10083) );
  INVX2TS U10240 ( .A(sa13[0]), .Y(n9859) );
  INVX2TS U10241 ( .A(sa00[2]), .Y(n9787) );
  INVX2TS U10242 ( .A(sa21[7]), .Y(n10330) );
  INVX2TS U10243 ( .A(sa13[5]), .Y(n9871) );
  INVX2TS U10244 ( .A(sa31[7]), .Y(n9373) );
  INVX2TS U10245 ( .A(sa13[7]), .Y(n9875) );
  INVX2TS U10246 ( .A(sa01[2]), .Y(n9344) );
  INVX2TS U10247 ( .A(sa21[3]), .Y(n10059) );
  INVX2TS U10248 ( .A(sa22[1]), .Y(n10079) );
  INVX2TS U10249 ( .A(sa13[4]), .Y(n9867) );
  INVX2TS U10250 ( .A(sa12[6]), .Y(n10075) );
  INVX2TS U10251 ( .A(sa23[7]), .Y(n9544) );
  INVX2TS U10252 ( .A(sa13[2]), .Y(n9863) );
  INVX2TS U10253 ( .A(sa00[4]), .Y(n9277) );
  INVX2TS U10254 ( .A(sa22[4]), .Y(n9450) );
  INVX2TS U10255 ( .A(sa23[5]), .Y(n9540) );
  INVX2TS U10256 ( .A(sa30[5]), .Y(n9819) );
  INVX2TS U10257 ( .A(sa02[0]), .Y(n10344) );
  INVX2TS U10258 ( .A(sa30[0]), .Y(n9807) );
  INVX2TS U10259 ( .A(sa12[7]), .Y(n9442) );
  INVX2TS U10260 ( .A(sa03[5]), .Y(n9529) );
  INVX2TS U10261 ( .A(sa03[7]), .Y(n10095) );
  INVX2TS U10262 ( .A(sa03[0]), .Y(n10358) );
  INVX2TS U10263 ( .A(sa03[3]), .Y(n10363) );
  INVX2TS U10264 ( .A(sa03[6]), .Y(n9855) );
  INVX2TS U10265 ( .A(sa03[1]), .Y(n9521) );
  INVX2TS U10266 ( .A(sa03[2]), .Y(n10091) );
  INVX2TS U10267 ( .A(sa03[4]), .Y(n9525) );
  INVX2TS U10268 ( .A(sa32[5]), .Y(n9847) );
  INVX2TS U10269 ( .A(sa32[7]), .Y(n10087) );
  INVX2TS U10270 ( .A(sa32[3]), .Y(n10353) );
  INVX2TS U10271 ( .A(sa32[0]), .Y(n9461) );
  INVX2TS U10272 ( .A(sa32[2]), .Y(n10348) );
  INVX2TS U10273 ( .A(sa32[4]), .Y(n9843) );
  INVX2TS U10274 ( .A(sa32[6]), .Y(n9851) );
  INVX2TS U10275 ( .A(sa20[2]), .Y(n10035) );
  INVX2TS U10276 ( .A(sa20[4]), .Y(n9795) );
  INVX2TS U10277 ( .A(sa20[6]), .Y(n10039) );
  INVX2TS U10278 ( .A(sa20[1]), .Y(n9285) );
  INVX2TS U10279 ( .A(sa20[0]), .Y(n9791) );
  INVX2TS U10280 ( .A(sa20[5]), .Y(n9799) );
  INVX2TS U10281 ( .A(sa20[7]), .Y(n9803) );
  INVX2TS U10282 ( .A(sa22[0]), .Y(n9839) );
  INVX2TS U10283 ( .A(n9381), .Y(n9383) );
  INVX2TS U10284 ( .A(n9488), .Y(n9490) );
  CLKBUFX2TS U10285 ( .A(n9041), .Y(n12655) );
  INVXLTS U10286 ( .A(w0[12]), .Y(n9314) );
  INVXLTS U10287 ( .A(w3[30]), .Y(n9614) );
  INVXLTS U10288 ( .A(w2[9]), .Y(n9478) );
  INVXLTS U10289 ( .A(w0[27]), .Y(n9336) );
  INVXLTS U10290 ( .A(w0[17]), .Y(n9319) );
  INVX2TS U10291 ( .A(n6927), .Y(n9793) );
  INVX2TS U10292 ( .A(n6927), .Y(n9794) );
  INVX1TS U10293 ( .A(n5197), .Y(n9276) );
  AOI22X1TS U10294 ( .A0(n6984), .A1(n9455), .B0(n6953), .B1(n1567), .Y(n7027)
         );
  INVX2TS U10295 ( .A(n6950), .Y(n9455) );
  INVX2TS U10296 ( .A(n5125), .Y(n9259) );
  AOI22X1TS U10297 ( .A0(n1358), .A1(n1407), .B0(n1408), .B1(n9777), .Y(n1406)
         );
  INVX2TS U10298 ( .A(n5147), .Y(n9267) );
  CLKINVX2TS U10299 ( .A(n1316), .Y(n9270) );
  INVX2TS U10300 ( .A(n1316), .Y(n9269) );
  CLKINVX2TS U10301 ( .A(n6950), .Y(n9456) );
  INVX2TS U10302 ( .A(n3331), .Y(n9073) );
  CLKINVX2TS U10303 ( .A(n5824), .Y(n9317) );
  CLKINVX2TS U10304 ( .A(n4024), .Y(n9125) );
  INVX1TS U10305 ( .A(n6991), .Y(n9460) );
  INVX1TS U10306 ( .A(n3381), .Y(n9088) );
  INVX1TS U10307 ( .A(n3381), .Y(n9089) );
  CLKINVX2TS U10308 ( .A(n2230), .Y(n9082) );
  INVX1TS U10309 ( .A(n3345), .Y(n9078) );
  INVX1TS U10310 ( .A(n3356), .Y(n9080) );
  CLKINVX2TS U10311 ( .A(n3356), .Y(n9081) );
  INVX1TS U10312 ( .A(n5824), .Y(n9318) );
  INVX2TS U10313 ( .A(n1361), .Y(n9776) );
  OAI22X1TS U10314 ( .A0(n9198), .A1(n1582), .B0(n9280), .B1(n5238), .Y(n5126)
         );
  OAI22X1TS U10315 ( .A0(n9184), .A1(n1596), .B0(n9093), .B1(n3441), .Y(n3332)
         );
  INVX2TS U10316 ( .A(n1529), .Y(n9212) );
  INVX1TS U10317 ( .A(n1402), .Y(n9235) );
  INVX2TS U10318 ( .A(n1294), .Y(n9783) );
  INVX1TS U10319 ( .A(n5157), .Y(n1770) );
  INVX1TS U10320 ( .A(n5174), .Y(n1647) );
  INVX2TS U10321 ( .A(n9752), .Y(n9753) );
  INVX2TS U10322 ( .A(n9202), .Y(n9203) );
  INVX1TS U10323 ( .A(n3420), .Y(n12657) );
  INVX2TS U10324 ( .A(n1481), .Y(n9227) );
  INVX1TS U10325 ( .A(n6932), .Y(n1644) );
  INVX1TS U10326 ( .A(n1340), .Y(n9255) );
  INVX1TS U10327 ( .A(n1384), .Y(n9243) );
  INVX1TS U10328 ( .A(n1481), .Y(n9228) );
  INVX2TS U10329 ( .A(n9273), .Y(n9274) );
  INVX1TS U10330 ( .A(n3363), .Y(n1784) );
  INVX2TS U10331 ( .A(n1384), .Y(n9242) );
  INVX2TS U10332 ( .A(n3380), .Y(n9085) );
  INVX2TS U10333 ( .A(n3380), .Y(n9084) );
  INVX2TS U10334 ( .A(n9223), .Y(n9224) );
  OAI22X1TS U10335 ( .A0(n1568), .A1(n6925), .B0(n9152), .B1(n7023), .Y(n6999)
         );
  INVX1TS U10336 ( .A(n1374), .Y(n9247) );
  INVX2TS U10337 ( .A(n9167), .Y(n9168) );
  INVX1TS U10338 ( .A(n1327), .Y(n9262) );
  INVX2TS U10339 ( .A(n9139), .Y(n9140) );
  INVX2TS U10340 ( .A(n1340), .Y(n9254) );
  INVX1TS U10341 ( .A(n3379), .Y(n1780) );
  INVX2TS U10342 ( .A(n5233), .Y(n9279) );
  INVX2TS U10343 ( .A(n9173), .Y(n9174) );
  INVX2TS U10344 ( .A(n5175), .Y(n9271) );
  INVX2TS U10345 ( .A(n1520), .Y(n9216) );
  INVX1TS U10346 ( .A(n1520), .Y(n9217) );
  INVX2TS U10347 ( .A(n1327), .Y(n9261) );
  INVX2TS U10348 ( .A(n3436), .Y(n9092) );
  INVX2TS U10349 ( .A(n1374), .Y(n9246) );
  INVX2TS U10350 ( .A(n1997), .Y(n9736) );
  INVX2TS U10351 ( .A(n5175), .Y(n9272) );
  INVX1TS U10352 ( .A(n1594), .Y(n10023) );
  INVX1TS U10353 ( .A(n3337), .Y(n1996) );
  INVX2TS U10354 ( .A(n1637), .Y(n10019) );
  INVX1TS U10355 ( .A(n5196), .Y(n1580) );
  INVX2TS U10356 ( .A(n1550), .Y(n9191) );
  INVX1TS U10357 ( .A(n1550), .Y(n9192) );
  INVXLTS U10358 ( .A(n6960), .Y(n12656) );
  INVX1TS U10359 ( .A(n1399), .Y(n1401) );
  INVX2TS U10360 ( .A(n1387), .Y(n9238) );
  INVX1TS U10361 ( .A(n9159), .Y(n9160) );
  INVX2TS U10362 ( .A(n1318), .Y(n9265) );
  INVX1TS U10363 ( .A(n9250), .Y(n9251) );
  INVX2TS U10364 ( .A(n1623), .Y(n9145) );
  INVX2TS U10365 ( .A(n1581), .Y(n9170) );
  INVX1TS U10366 ( .A(n1318), .Y(n9266) );
  INVX2TS U10367 ( .A(n1595), .Y(n9163) );
  INVX2TS U10368 ( .A(n1474), .Y(n9230) );
  INVX1TS U10369 ( .A(n1474), .Y(n9231) );
  INVX2TS U10370 ( .A(n1305), .Y(n9779) );
  CLKINVX2TS U10371 ( .A(n9136), .Y(n9137) );
  CLKINVX2TS U10372 ( .A(n1597), .Y(n9159) );
  INVX2TS U10373 ( .A(n1557), .Y(n9181) );
  CLKINVX2TS U10374 ( .A(n9148), .Y(n9149) );
  INVX1TS U10375 ( .A(n1557), .Y(n9182) );
  INVX1TS U10376 ( .A(n7023), .Y(n1568) );
  INVX1TS U10377 ( .A(n6990), .Y(n1566) );
  INVX1TS U10378 ( .A(n1395), .Y(n1398) );
  AOI211X1TS U10379 ( .A0(n11781), .A1(n9098), .B0(n3637), .C0(n3638), .Y(
        n3634) );
  AOI211X1TS U10380 ( .A0(n12248), .A1(n12409), .B0(n5884), .C0(n5885), .Y(
        n5883) );
  AOI211X1TS U10381 ( .A0(n12260), .A1(n12437), .B0(n4028), .C0(n4029), .Y(
        n4027) );
  AOI211X1TS U10382 ( .A0(n11283), .A1(n11699), .B0(n6825), .C0(n6826), .Y(
        n6824) );
  AOI211X1TS U10383 ( .A0(n11233), .A1(n11681), .B0(n6767), .C0(n6768), .Y(
        n6766) );
  AOI211X1TS U10384 ( .A0(n12237), .A1(n12421), .B0(n4084), .C0(n4085), .Y(
        n4083) );
  AOI211X1TS U10385 ( .A0(n11368), .A1(n11750), .B0(n4968), .C0(n4969), .Y(
        n4967) );
  AOI211X1TS U10386 ( .A0(n12225), .A1(n12393), .B0(n5828), .C0(n5829), .Y(
        n5827) );
  AOI211X1TS U10387 ( .A0(n11320), .A1(n11731), .B0(n5026), .C0(n5027), .Y(
        n5025) );
  OAI32X1TS U10388 ( .A0(n7160), .A1(n12107), .A2(n12551), .B0(n11462), .B1(
        n7160), .Y(n7084) );
  AOI211X1TS U10389 ( .A0(n10549), .A1(n12279), .B0(n6291), .C0(n6292), .Y(
        n6290) );
  AOI211X1TS U10390 ( .A0(n12487), .A1(n12363), .B0(n8013), .C0(n8014), .Y(
        n8012) );
  AOI211X1TS U10391 ( .A0(n12518), .A1(n6133), .B0(n6494), .C0(n6838), .Y(
        n6823) );
  AOI211X1TS U10392 ( .A0(n11327), .A1(n12436), .B0(n4148), .C0(n4149), .Y(
        n4146) );
  AOI211X1TS U10393 ( .A0(n12506), .A1(n4223), .B0(n4694), .C0(n5039), .Y(
        n5024) );
  AOI211X1TS U10394 ( .A0(n11809), .A1(n12378), .B0(n4787), .C0(n4788), .Y(
        n4786) );
  AOI22X1TS U10395 ( .A0(n11544), .A1(n12341), .B0(n12454), .B1(n9094), .Y(
        n3033) );
  AOI211X1TS U10396 ( .A0(n12523), .A1(n4179), .B0(n4622), .C0(n4981), .Y(
        n4966) );
  AOI211X1TS U10397 ( .A0(n11276), .A1(n12392), .B0(n6058), .C0(n6059), .Y(
        n6056) );
  AOI211X1TS U10398 ( .A0(n11324), .A1(n12408), .B0(n6102), .C0(n6103), .Y(
        n6100) );
  AOI211X1TS U10399 ( .A0(n11812), .A1(n8162), .B0(n7950), .C0(n8163), .Y(
        n7371) );
  AOI211X1TS U10400 ( .A0(n12503), .A1(n6089), .B0(n6422), .C0(n6780), .Y(
        n6765) );
  AOI211X1TS U10401 ( .A0(n11279), .A1(n12420), .B0(n4192), .C0(n4193), .Y(
        n4190) );
  AOI211X1TS U10402 ( .A0(n11980), .A1(n12450), .B0(n6587), .C0(n6588), .Y(
        n6586) );
  AOI22X1TS U10403 ( .A0(n12526), .A1(n9372), .B0(n11710), .B1(n12274), .Y(
        n6501) );
  AOI211X1TS U10404 ( .A0(n11123), .A1(n12487), .B0(n7740), .C0(n8329), .Y(
        n7634) );
  AOI22X1TS U10405 ( .A0(n12448), .A1(n5784), .B0(n12574), .B1(n6183), .Y(
        n6182) );
  AOI22X1TS U10406 ( .A0(n12500), .A1(n9166), .B0(n11721), .B1(n12215), .Y(
        n4701) );
  AOI22X1TS U10407 ( .A0(n11758), .A1(n9353), .B0(n12536), .B1(n6289), .Y(
        n6283) );
  AOI22X1TS U10408 ( .A0(n11739), .A1(n9157), .B0(n11751), .B1(n4414), .Y(
        n4410) );
  AOI22X1TS U10409 ( .A0(n11712), .A1(n9371), .B0(n11699), .B1(n6257), .Y(
        n6253) );
  AOI211X1TS U10410 ( .A0(n3924), .A1(n9099), .B0(n4472), .C0(n4473), .Y(n4470) );
  AOI22X1TS U10411 ( .A0(n10952), .A1(n5784), .B0(n9637), .B1(n6027), .Y(n6021) );
  AOI22X1TS U10412 ( .A0(n10800), .A1(n3990), .B0(n9634), .B1(n4260), .Y(n4253) );
  AOI22X1TS U10413 ( .A0(n12517), .A1(n9158), .B0(n11737), .B1(n12222), .Y(
        n4629) );
  AOI22X1TS U10414 ( .A0(n12510), .A1(n9364), .B0(n11692), .B1(n12266), .Y(
        n6429) );
  AOI22X1TS U10415 ( .A0(n11676), .A1(n5783), .B0(n9637), .B1(n5784), .Y(n5776) );
  OAI2BB2XLTS U10416 ( .B0(n6341), .B1(n12285), .A0N(n6372), .A1N(n11759), .Y(
        n6869) );
  OAI32X1TS U10417 ( .A0(n11441), .A1(n3024), .A2(n11816), .B0(n11829), .B1(
        n3024), .Y(n3023) );
  INVX2TS U10418 ( .A(n2057), .Y(n9094) );
  AOI22X1TS U10419 ( .A0(n11694), .A1(n9363), .B0(n11682), .B1(n6217), .Y(
        n6213) );
  AOI22X1TS U10420 ( .A0(n11720), .A1(n9165), .B0(n11733), .B1(n4454), .Y(
        n4450) );
  AOI22X1TS U10421 ( .A0(n11787), .A1(n3989), .B0(n12594), .B1(n3990), .Y(
        n3988) );
  AOI22X1TS U10422 ( .A0(n12376), .A1(n3990), .B0(n12592), .B1(n4379), .Y(
        n4378) );
  AOI221X1TS U10423 ( .A0(n11543), .A1(n2665), .B0(n12651), .B1(n2491), .C0(
        n2666), .Y(n2664) );
  CLKINVX2TS U10424 ( .A(n7335), .Y(n9492) );
  AOI211X1TS U10425 ( .A0(n11974), .A1(n12512), .B0(n5879), .C0(n6756), .Y(
        n6075) );
  AOI221X1TS U10426 ( .A0(n11768), .A1(n10390), .B0(n12016), .B1(n4837), .C0(
        n4873), .Y(n4872) );
  AOI211X1TS U10427 ( .A0(n12511), .A1(n10581), .B0(n6406), .C0(n6794), .Y(
        n6077) );
  OAI31X1TS U10428 ( .A0(n9903), .A1(n11792), .A2(n9095), .B0(n9634), .Y(n4233) );
  AOI211X1TS U10429 ( .A0(n11680), .A1(n12235), .B0(n5454), .C0(n5455), .Y(
        n5452) );
  CLKINVX2TS U10430 ( .A(n7364), .Y(n9829) );
  AOI211X1TS U10431 ( .A0(n12232), .A1(n6426), .B0(n6757), .C0(n6758), .Y(
        n6074) );
  INVX2TS U10432 ( .A(n7459), .Y(n9515) );
  AOI211X1TS U10433 ( .A0(n12255), .A1(n6498), .B0(n6815), .C0(n6816), .Y(
        n6118) );
  AOI211X1TS U10434 ( .A0(n11971), .A1(n12528), .B0(n5935), .C0(n6814), .Y(
        n6119) );
  AOI211X1TS U10435 ( .A0(n12621), .A1(n3924), .B0(n4867), .C0(n4497), .Y(
        n4861) );
  AOI22X1TS U10436 ( .A0(n9903), .A1(n12046), .B0(n10881), .B1(n11786), .Y(
        n3623) );
  AOI211X1TS U10437 ( .A0(n11698), .A1(n12258), .B0(n5520), .C0(n5521), .Y(
        n5518) );
  AOI22X1TS U10438 ( .A0(n10434), .A1(n10430), .B0(n12074), .B1(n12043), .Y(
        n3828) );
  AOI211X1TS U10439 ( .A0(n12228), .A1(n4698), .B0(n5016), .C0(n5017), .Y(
        n4208) );
  INVX2TS U10440 ( .A(n1823), .Y(n9748) );
  AOI21X1TS U10441 ( .A0(n12500), .A1(n12509), .B0(n5041), .Y(n4210) );
  AOI211X1TS U10442 ( .A0(n12501), .A1(n10409), .B0(n4678), .C0(n5053), .Y(
        n4211) );
  AOI211X1TS U10443 ( .A0(n12517), .A1(n10404), .B0(n4606), .C0(n4995), .Y(
        n4167) );
  INVX1TS U10444 ( .A(n6070), .Y(n9364) );
  AOI22X1TS U10445 ( .A0(n11829), .A1(n10195), .B0(n12453), .B1(n2642), .Y(
        n2631) );
  AOI21X1TS U10446 ( .A0(n12514), .A1(n12522), .B0(n4983), .Y(n4166) );
  INVX2TS U10447 ( .A(n7335), .Y(n9491) );
  INVX2TS U10448 ( .A(n1823), .Y(n9749) );
  AOI21X1TS U10449 ( .A0(n12512), .A1(n12505), .B0(n6782), .Y(n6076) );
  INVX1TS U10450 ( .A(n8175), .Y(n9511) );
  AOI211X1TS U10451 ( .A0(n10248), .A1(n11841), .B0(n2455), .C0(n2818), .Y(
        n2817) );
  AOI211X1TS U10452 ( .A0(n12624), .A1(n12452), .B0(n3080), .C0(n3081), .Y(
        n3079) );
  INVX1TS U10453 ( .A(n4204), .Y(n9166) );
  AOI21X1TS U10454 ( .A0(n12529), .A1(n12518), .B0(n6840), .Y(n6120) );
  AOI211X1TS U10455 ( .A0(n12052), .A1(n12500), .B0(n4135), .C0(n5015), .Y(
        n4209) );
  AOI211X1TS U10456 ( .A0(n12251), .A1(n4626), .B0(n4958), .C0(n4959), .Y(
        n4164) );
  AOI21X1TS U10457 ( .A0(n10589), .A1(n12454), .B0(n3068), .Y(n3066) );
  OAI31X1TS U10458 ( .A0(n9954), .A1(n11678), .A2(n9284), .B0(n12576), .Y(
        n6000) );
  AOI211X1TS U10459 ( .A0(n12058), .A1(n12515), .B0(n4079), .C0(n4957), .Y(
        n4165) );
  AOI211X1TS U10460 ( .A0(n12046), .A1(n4260), .B0(n4754), .C0(n4772), .Y(
        n4937) );
  INVX1TS U10461 ( .A(n6114), .Y(n9372) );
  AOI211X1TS U10462 ( .A0(n11909), .A1(n12345), .B0(n8185), .C0(n8186), .Y(
        n8184) );
  INVX1TS U10463 ( .A(n5973), .Y(n9353) );
  INVX1TS U10464 ( .A(n4160), .Y(n9158) );
  AOI22X1TS U10465 ( .A0(n11135), .A1(n1844), .B0(n10972), .B1(n9760), .Y(
        n3161) );
  INVX2TS U10466 ( .A(n7121), .Y(n9805) );
  AOI221X1TS U10467 ( .A0(n11840), .A1(n1933), .B0(n11924), .B1(n12602), .C0(
        n2849), .Y(n1734) );
  AOI221X1TS U10468 ( .A0(n11846), .A1(n1870), .B0(n11936), .B1(n12598), .C0(
        n2925), .Y(n1696) );
  AOI211X1TS U10469 ( .A0(n11536), .A1(n12653), .B0(n3051), .C0(n3280), .Y(
        n3279) );
  AOI211X1TS U10470 ( .A0(n10195), .A1(n12289), .B0(n2779), .C0(n2780), .Y(
        n2778) );
  AOI211X1TS U10471 ( .A0(n12288), .A1(n11537), .B0(n3042), .C0(n2639), .Y(
        n3040) );
  INVX2TS U10472 ( .A(n7459), .Y(n9516) );
  CLKINVX2TS U10473 ( .A(n7121), .Y(n9806) );
  AOI211X1TS U10474 ( .A0(n12045), .A1(n4244), .B0(n4770), .C0(n4771), .Y(
        n4768) );
  INVX2TS U10475 ( .A(n7364), .Y(n9830) );
  AOI211X1TS U10476 ( .A0(n12526), .A1(n10585), .B0(n6478), .C0(n6852), .Y(
        n6121) );
  INVX2TS U10477 ( .A(n7359), .Y(n9825) );
  OAI32X1TS U10478 ( .A0(n5486), .A1(n12218), .A2(n12391), .B0(n9958), .B1(
        n5486), .Y(n5470) );
  AOI22X1TS U10479 ( .A0(n11542), .A1(n12105), .B0(n12651), .B1(n11009), .Y(
        n2155) );
  OAI32X1TS U10480 ( .A0(n5552), .A1(n12241), .A2(n12407), .B0(n9962), .B1(
        n5552), .Y(n5536) );
  OAI32X1TS U10481 ( .A0(n7968), .A1(n11086), .A2(n12345), .B0(n11499), .B1(
        n7968), .Y(n7965) );
  AOI211X1TS U10482 ( .A0(n11758), .A1(n12434), .B0(n6623), .C0(n6902), .Y(
        n5963) );
  CLKINVX1TS U10483 ( .A(n7339), .Y(n11866) );
  AOI22X1TS U10484 ( .A0(n11703), .A1(n4306), .B0(n12018), .B1(n4307), .Y(
        n4298) );
  AOI211X1TS U10485 ( .A0(n11452), .A1(n12326), .B0(n3006), .C0(n3007), .Y(
        n3005) );
  OAI32X1TS U10486 ( .A0(n3797), .A1(n12245), .A2(n12422), .B0(n9910), .B1(
        n3797), .Y(n3781) );
  INVX2TS U10487 ( .A(n1956), .Y(n9104) );
  INVX1TS U10488 ( .A(n2202), .Y(n9087) );
  INVX2TS U10489 ( .A(n6341), .Y(n9407) );
  INVX2TS U10490 ( .A(n12442), .Y(n9954) );
  INVX2TS U10491 ( .A(n5806), .Y(n9312) );
  CLKINVX2TS U10492 ( .A(n7315), .Y(n10652) );
  INVX2TS U10493 ( .A(n10791), .Y(n10116) );
  AOI211X1TS U10494 ( .A0(n12576), .A1(n9998), .B0(n6570), .C0(n6020), .Y(
        n6695) );
  CLKINVX2TS U10495 ( .A(n1956), .Y(n9105) );
  INVX2TS U10496 ( .A(n1728), .Y(n9761) );
  OAI31X1TS U10497 ( .A0(n12651), .A1(n12111), .A2(n12104), .B0(n12615), .Y(
        n3064) );
  OAI32X1TS U10498 ( .A0(n3731), .A1(n12268), .A2(n12435), .B0(n9906), .B1(
        n3731), .Y(n3715) );
  AOI211X1TS U10499 ( .A0(n12594), .A1(n10130), .B0(n4770), .C0(n4252), .Y(
        n4896) );
  AOI22X1TS U10500 ( .A0(n12488), .A1(n7330), .B0(n11592), .B1(n7825), .Y(
        n8025) );
  INVX2TS U10501 ( .A(n11373), .Y(n10238) );
  INVX1TS U10502 ( .A(n10983), .Y(n10491) );
  INVX2TS U10503 ( .A(n1766), .Y(n9756) );
  AOI22X1TS U10504 ( .A0(n11958), .A1(n7825), .B0(n12184), .B1(n7487), .Y(
        n8331) );
  CLKINVX1TS U10505 ( .A(n5806), .Y(n9313) );
  OAI31X1TS U10506 ( .A0(n12291), .A1(n12653), .A2(n10183), .B0(n11028), .Y(
        n3078) );
  AOI22X1TS U10507 ( .A0(n11856), .A1(n11958), .B0(n12371), .B1(n7487), .Y(
        n8445) );
  AOI221X1TS U10508 ( .A0(n11828), .A1(n12311), .B0(n12453), .B1(n12106), .C0(
        n3283), .Y(n3282) );
  AOI22X1TS U10509 ( .A0(n12652), .A1(n2070), .B0(n10183), .B1(n11068), .Y(
        n3025) );
  INVX2TS U10510 ( .A(n12390), .Y(n9904) );
  CLKINVX2TS U10511 ( .A(n10668), .Y(n10010) );
  AOI211X1TS U10512 ( .A0(n12071), .A1(n12377), .B0(n4778), .C0(n4891), .Y(
        n4890) );
  AOI22X1TS U10513 ( .A0(n10179), .A1(n11502), .B0(n11520), .B1(n2549), .Y(
        n3090) );
  AOI211X1TS U10514 ( .A0(n11791), .A1(n12376), .B0(n3816), .C0(n4269), .Y(
        n4267) );
  INVX2TS U10515 ( .A(n12439), .Y(n9953) );
  INVX2TS U10516 ( .A(n11372), .Y(n10237) );
  INVX2TS U10517 ( .A(n10791), .Y(n10115) );
  AOI22X1TS U10518 ( .A0(n10516), .A1(n11442), .B0(n12104), .B1(n9689), .Y(
        n3277) );
  INVX2TS U10519 ( .A(n1766), .Y(n9757) );
  AOI211X1TS U10520 ( .A0(n12391), .A1(n12227), .B0(n6745), .C0(n6746), .Y(
        n6744) );
  INVX2TS U10521 ( .A(n10984), .Y(n10492) );
  INVX1TS U10522 ( .A(n11019), .Y(n10193) );
  INVX2TS U10523 ( .A(n7067), .Y(n9797) );
  CLKINVX2TS U10524 ( .A(n4303), .Y(n9938) );
  INVX2TS U10525 ( .A(n5658), .Y(n10969) );
  INVX2TS U10526 ( .A(n5658), .Y(n10968) );
  AOI21X1TS U10527 ( .A0(n11206), .A1(n5296), .B0(n6597), .Y(n6595) );
  OAI21X1TS U10528 ( .A0(n10168), .A1(n11501), .B0(n11518), .Y(n3088) );
  AOI211X1TS U10529 ( .A0(n12435), .A1(n12262), .B0(n4946), .C0(n4947), .Y(
        n4945) );
  INVX2TS U10530 ( .A(n12387), .Y(n9903) );
  INVX2TS U10531 ( .A(n10668), .Y(n10009) );
  AOI22X1TS U10532 ( .A0(n11267), .A1(n10121), .B0(n12043), .B1(n3822), .Y(
        n4790) );
  CLKINVX2TS U10533 ( .A(n7339), .Y(n11867) );
  AOI211X1TS U10534 ( .A0(n11845), .A1(n3163), .B0(n1866), .C0(n3164), .Y(
        n3162) );
  CLKINVX2TS U10535 ( .A(n4303), .Y(n9937) );
  INVX2TS U10536 ( .A(n2202), .Y(n9086) );
  INVX1TS U10537 ( .A(n10757), .Y(n10433) );
  INVX2TS U10538 ( .A(n1728), .Y(n9760) );
  AOI211X1TS U10539 ( .A0(n12324), .A1(n12647), .B0(n2954), .C0(n2955), .Y(
        n2181) );
  AOI22X1TS U10540 ( .A0(n10515), .A1(n3031), .B0(n12453), .B1(n12106), .Y(
        n3030) );
  INVX2TS U10541 ( .A(n10758), .Y(n10434) );
  INVX2TS U10542 ( .A(n7339), .Y(n11868) );
  INVX2TS U10543 ( .A(n3504), .Y(n9096) );
  INVX2TS U10544 ( .A(n3917), .Y(n9118) );
  INVX2TS U10545 ( .A(n7209), .Y(n9813) );
  OAI31X1TS U10546 ( .A0(n11677), .A1(n5316), .A2(n6162), .B0(n9375), .Y(n6166) );
  INVX2TS U10547 ( .A(n4020), .Y(n9121) );
  AOI211X1TS U10548 ( .A0(n12594), .A1(n11811), .B0(n4754), .C0(n3981), .Y(
        n4753) );
  AOI21X1TS U10549 ( .A0(n11416), .A1(n3498), .B0(n4797), .Y(n4795) );
  OAI31X1TS U10550 ( .A0(n11560), .A1(n12338), .A2(n12650), .B0(n12451), .Y(
        n1966) );
  INVX2TS U10551 ( .A(n11019), .Y(n10194) );
  INVX2TS U10552 ( .A(n3504), .Y(n9095) );
  OAI31X1TS U10553 ( .A0(n11791), .A1(n3518), .A2(n4358), .B0(n9179), .Y(n4362) );
  CLKINVX2TS U10554 ( .A(n7698), .Y(n9858) );
  INVX1TS U10555 ( .A(n5658), .Y(n10970) );
  INVX1TS U10556 ( .A(n1668), .Y(n12187) );
  CLKINVX2TS U10557 ( .A(n11329), .Y(n9388) );
  INVX2TS U10558 ( .A(n10899), .Y(n11302) );
  INVX2TS U10559 ( .A(n10780), .Y(n11315) );
  AOI22X1TS U10560 ( .A0(n11738), .A1(n4964), .B0(n9647), .B1(n3542), .Y(n4962) );
  AOI22X1TS U10561 ( .A0(n4203), .A1(n11719), .B0(n11280), .B1(n3581), .Y(
        n4123) );
  CLKINVX2TS U10562 ( .A(n3984), .Y(n10107) );
  AOI221X1TS U10563 ( .A0(n11929), .A1(n11131), .B0(n12365), .B1(n12603), .C0(
        n1748), .Y(n1742) );
  AOI211X1TS U10564 ( .A0(n9647), .A1(n12251), .B0(n3856), .C0(n4071), .Y(
        n4070) );
  OAI2BB2XLTS U10565 ( .B0(n6460), .B1(n10919), .A0N(n5540), .A1N(n12258), .Y(
        n6808) );
  INVX2TS U10566 ( .A(n5548), .Y(n9307) );
  INVX2TS U10567 ( .A(n12419), .Y(n10131) );
  CLKINVX2TS U10568 ( .A(n11002), .Y(n11239) );
  AOI211X1TS U10569 ( .A0(n10913), .A1(n11281), .B0(n5509), .C0(n5510), .Y(
        n5504) );
  AOI22X1TS U10570 ( .A0(n12511), .A1(n10458), .B0(n11688), .B1(n12036), .Y(
        n6207) );
  INVX1TS U10571 ( .A(n1689), .Y(n10680) );
  CLKINVX2TS U10572 ( .A(n10779), .Y(n11316) );
  INVX2TS U10573 ( .A(n10852), .Y(n11252) );
  INVX2TS U10574 ( .A(n12394), .Y(n10158) );
  AOI22X1TS U10575 ( .A0(n12436), .A1(n11356), .B0(n12587), .B1(n11737), .Y(
        n4996) );
  INVX2TS U10576 ( .A(n3636), .Y(n9098) );
  OAI31X1TS U10577 ( .A0(n12370), .A1(n12487), .A2(n12141), .B0(n12189), .Y(
        n8450) );
  AOI22X1TS U10578 ( .A0(n11847), .A1(n2701), .B0(n10972), .B1(n2093), .Y(
        n2693) );
  INVX1TS U10579 ( .A(n5482), .Y(n9298) );
  INVX2TS U10580 ( .A(n12216), .Y(n9663) );
  AOI211X1TS U10581 ( .A0(n12576), .A1(n11980), .B0(n6554), .C0(n5813), .Y(
        n6553) );
  AOI22X1TS U10582 ( .A0(n11693), .A1(n6763), .B0(n9730), .B1(n5340), .Y(n6761) );
  INVX1TS U10583 ( .A(n3793), .Y(n9115) );
  CLKINVX2TS U10584 ( .A(n9190), .Y(n12207) );
  OAI2BB2XLTS U10585 ( .B0(n6388), .B1(n10891), .A0N(n5474), .A1N(n12235), .Y(
        n6750) );
  INVX1TS U10586 ( .A(n10853), .Y(n11253) );
  INVX2TS U10587 ( .A(n12391), .Y(n10157) );
  INVX2TS U10588 ( .A(n12438), .Y(n10140) );
  AOI22X1TS U10589 ( .A0(n12527), .A1(n10466), .B0(n11706), .B1(n12050), .Y(
        n6247) );
  AOI22X1TS U10590 ( .A0(n10270), .A1(n12456), .B0(n11813), .B1(n12552), .Y(
        n7152) );
  OAI31X1TS U10591 ( .A0(n11885), .A1(n11814), .A2(n11431), .B0(n12551), .Y(
        n7804) );
  CLKINVX2TS U10592 ( .A(n10869), .Y(n11301) );
  INVX2TS U10593 ( .A(n5797), .Y(n10206) );
  CLKINVX2TS U10594 ( .A(n9189), .Y(n12206) );
  AOI221X1TS U10595 ( .A0(n11943), .A1(n11152), .B0(n12374), .B1(n12600), .C0(
        n1710), .Y(n1704) );
  CLKINVX2TS U10596 ( .A(n5797), .Y(n10205) );
  INVX2TS U10597 ( .A(n10954), .Y(n11500) );
  AOI22X1TS U10598 ( .A0(n12499), .A1(n10442), .B0(n11726), .B1(n11988), .Y(
        n4444) );
  CLKINVX2TS U10599 ( .A(n11001), .Y(n11240) );
  AOI22X1TS U10600 ( .A0(n12220), .A1(n11692), .B0(n11275), .B1(n5340), .Y(
        n5867) );
  CLKINVX2TS U10601 ( .A(n10900), .Y(n11304) );
  AOI211X1TS U10602 ( .A0(n9731), .A1(n12232), .B0(n5686), .C0(n5871), .Y(
        n5870) );
  CLKINVX2TS U10603 ( .A(n11000), .Y(n11241) );
  INVX2TS U10604 ( .A(n12265), .Y(n9702) );
  AOI22X1TS U10605 ( .A0(n11957), .A1(n11551), .B0(n11898), .B1(n11860), .Y(
        n8293) );
  AOI22X1TS U10606 ( .A0(n12267), .A1(n11738), .B0(n11327), .B1(n3542), .Y(
        n4067) );
  INVX2TS U10607 ( .A(n10956), .Y(n11501) );
  CLKINVX2TS U10608 ( .A(n11022), .Y(n11079) );
  AOI22X1TS U10609 ( .A0(n12063), .A1(n6633), .B0(n12281), .B1(n9978), .Y(
        n6621) );
  AOI211X1TS U10610 ( .A0(n10885), .A1(n11235), .B0(n5443), .C0(n5444), .Y(
        n5438) );
  AOI22X1TS U10611 ( .A0(n11246), .A1(n9635), .B0(n12224), .B1(n12233), .Y(
        n6743) );
  AOI22X1TS U10612 ( .A0(n12392), .A1(n11247), .B0(n5875), .B1(n11693), .Y(
        n6795) );
  INVX1TS U10613 ( .A(n10915), .Y(n11352) );
  AOI22X1TS U10614 ( .A0(n11856), .A1(n7826), .B0(n11552), .B1(n12486), .Y(
        n8426) );
  INVX2TS U10615 ( .A(n5482), .Y(n9297) );
  INVX2TS U10616 ( .A(n2033), .Y(n11051) );
  INVX2TS U10617 ( .A(n3984), .Y(n10108) );
  INVX2TS U10618 ( .A(n3727), .Y(n9106) );
  CLKINVX2TS U10619 ( .A(n9990), .Y(n10830) );
  INVX2TS U10620 ( .A(n5302), .Y(n9283) );
  INVX2TS U10621 ( .A(n3793), .Y(n9114) );
  AOI22X1TS U10622 ( .A0(n11508), .A1(n11519), .B0(n11954), .B1(n12182), .Y(
        n2967) );
  AOI22X1TS U10623 ( .A0(n12420), .A1(n11310), .B0(n12579), .B1(n11720), .Y(
        n5054) );
  AOI22X1TS U10624 ( .A0(n12408), .A1(n11293), .B0(n12591), .B1(n11710), .Y(
        n6853) );
  AOI22X1TS U10625 ( .A0(n11208), .A1(n5808), .B0(n11668), .B1(n6046), .Y(
        n6044) );
  CLKINVX2TS U10626 ( .A(n3668), .Y(n9670) );
  INVX2TS U10627 ( .A(n7608), .Y(n9531) );
  INVX2TS U10628 ( .A(n12435), .Y(n10139) );
  INVX2TS U10629 ( .A(n10597), .Y(n10183) );
  AOI22X1TS U10630 ( .A0(n11416), .A1(n4022), .B0(n12044), .B1(n4279), .Y(
        n4277) );
  OAI2BB2XLTS U10631 ( .B0(n11576), .B1(n12129), .A0N(n8219), .A1N(n12342), 
        .Y(n8218) );
  INVX2TS U10632 ( .A(n1668), .Y(n12186) );
  CLKINVX2TS U10633 ( .A(n10768), .Y(n11363) );
  AOI22X1TS U10634 ( .A0(n10081), .A1(n11516), .B0(n12486), .B1(n10316), .Y(
        n8281) );
  CLKINVX2TS U10635 ( .A(n11012), .Y(n11288) );
  INVX1TS U10636 ( .A(n5548), .Y(n9308) );
  CLKINVX2TS U10637 ( .A(n9934), .Y(n10939) );
  AOI221X1TS U10638 ( .A0(n12650), .A1(n10519), .B0(n12613), .B1(n10949), .C0(
        n3032), .Y(n3028) );
  OAI2BB2XLTS U10639 ( .B0(n4660), .B1(n10821), .A0N(n3785), .A1N(n12230), .Y(
        n5009) );
  AOI22X1TS U10640 ( .A0(n10805), .A1(n11733), .B0(n11308), .B1(n12228), .Y(
        n4666) );
  AOI22X1TS U10641 ( .A0(n12240), .A1(n11711), .B0(n11324), .B1(n5379), .Y(
        n5923) );
  AOI22X1TS U10642 ( .A0(n11357), .A1(n9636), .B0(n12259), .B1(n12252), .Y(
        n4944) );
  INVX2TS U10643 ( .A(n10916), .Y(n11351) );
  CLKINVX2TS U10644 ( .A(n3701), .Y(n9667) );
  INVX1TS U10645 ( .A(n10619), .Y(n12105) );
  INVX1TS U10646 ( .A(n3727), .Y(n9107) );
  INVX1TS U10647 ( .A(n5302), .Y(n9284) );
  AOI211X1TS U10648 ( .A0(n9735), .A1(n12255), .B0(n5711), .C0(n5927), .Y(
        n5926) );
  CLKINVX2TS U10649 ( .A(n11023), .Y(n11081) );
  AOI22X1TS U10650 ( .A0(n10908), .A1(n11682), .B0(n11245), .B1(n12233), .Y(
        n6394) );
  CLKINVX2TS U10651 ( .A(n1986), .Y(n11554) );
  AOI22X1TS U10652 ( .A0(n11711), .A1(n6821), .B0(n9735), .B1(n5379), .Y(n6819) );
  CLKINVX2TS U10653 ( .A(n10589), .Y(n11550) );
  INVX2TS U10654 ( .A(n1968), .Y(n11560) );
  AOI22X1TS U10655 ( .A0(n12515), .A1(n10451), .B0(n11744), .B1(n12003), .Y(
        n4404) );
  INVX1TS U10656 ( .A(n1689), .Y(n10679) );
  CLKINVX2TS U10657 ( .A(n10778), .Y(n11314) );
  AOI211X1TS U10658 ( .A0(n10674), .A1(n11813), .B0(n7423), .C0(n7424), .Y(
        n7420) );
  INVX2TS U10659 ( .A(n12422), .Y(n10132) );
  CLKINVX2TS U10660 ( .A(n11013), .Y(n11289) );
  AOI22X1TS U10661 ( .A0(n10701), .A1(n11505), .B0(n12344), .B1(n11497), .Y(
        n8214) );
  AOI22X1TS U10662 ( .A0(n10831), .A1(n11749), .B0(n11357), .B1(n12252), .Y(
        n4594) );
  AOI22X1TS U10663 ( .A0(n11956), .A1(n12190), .B0(n11096), .B1(n11146), .Y(
        n8330) );
  INVX2TS U10664 ( .A(n7608), .Y(n9532) );
  CLKINVX2TS U10665 ( .A(n10767), .Y(n11364) );
  INVX1TS U10666 ( .A(n10955), .Y(n11502) );
  AOI22X1TS U10667 ( .A0(n11719), .A1(n5022), .B0(n9642), .B1(n3581), .Y(n5020) );
  AOI22X1TS U10668 ( .A0(n10917), .A1(n4179), .B0(n10906), .B1(n12253), .Y(
        n4172) );
  AOI211X1TS U10669 ( .A0(n10556), .A1(n12368), .B0(n2827), .C0(n2828), .Y(
        n2825) );
  INVX2TS U10670 ( .A(n2033), .Y(n11052) );
  AOI22X1TS U10671 ( .A0(n12605), .A1(n11132), .B0(n11841), .B1(n2719), .Y(
        n2824) );
  OAI2BB2XLTS U10672 ( .B0(n4588), .B1(n10849), .A0N(n3719), .A1N(n12254), .Y(
        n4951) );
  INVX2TS U10673 ( .A(n12410), .Y(n10166) );
  CLKINVX2TS U10674 ( .A(n10901), .Y(n11303) );
  OAI21X1TS U10675 ( .A0(n11551), .A1(n11098), .B0(n12488), .Y(n7661) );
  AOI22X1TS U10676 ( .A0(n12646), .A1(n11424), .B0(n12195), .B1(n12180), .Y(
        n2950) );
  AOI22X1TS U10677 ( .A0(n11827), .A1(n2657), .B0(n11817), .B1(n12290), .Y(
        n3050) );
  AOI22X1TS U10678 ( .A0(n10870), .A1(n6133), .B0(n10879), .B1(n12257), .Y(
        n6126) );
  AOI22X1TS U10679 ( .A0(n11768), .A1(n10133), .B0(n9189), .B1(n12016), .Y(
        n4490) );
  INVX2TS U10680 ( .A(n1968), .Y(n11562) );
  INVX2TS U10681 ( .A(n10597), .Y(n10184) );
  INVX2TS U10682 ( .A(n3701), .Y(n9666) );
  INVX2TS U10683 ( .A(n3636), .Y(n9099) );
  INVX2TS U10684 ( .A(n12215), .Y(n9662) );
  AOI22X1TS U10685 ( .A0(n12339), .A1(n3058), .B0(n12289), .B1(n12310), .Y(
        n3054) );
  AOI22X1TS U10686 ( .A0(n10935), .A1(n11700), .B0(n11294), .B1(n12256), .Y(
        n6466) );
  INVX2TS U10687 ( .A(n1968), .Y(n11561) );
  INVX2TS U10688 ( .A(n10621), .Y(n12104) );
  INVX2TS U10689 ( .A(n12407), .Y(n10165) );
  CLKINVX2TS U10690 ( .A(n10766), .Y(n11362) );
  INVX2TS U10691 ( .A(n10620), .Y(n12106) );
  AOI22X1TS U10692 ( .A0(n11840), .A1(n2734), .B0(n10988), .B1(n2119), .Y(
        n2726) );
  CLKINVX2TS U10693 ( .A(n2628), .Y(n10508) );
  CLKINVX2TS U10694 ( .A(n1986), .Y(n11556) );
  INVX2TS U10695 ( .A(n12273), .Y(n9706) );
  INVX2TS U10696 ( .A(n12398), .Y(n9643) );
  INVX2TS U10697 ( .A(n10387), .Y(n11725) );
  AOI22X1TS U10698 ( .A0(n11822), .A1(n11452), .B0(n11514), .B1(n2577), .Y(
        n3113) );
  INVX1TS U10699 ( .A(n7651), .Y(n12363) );
  INVX2TS U10700 ( .A(n12398), .Y(n9642) );
  INVX2TS U10701 ( .A(n4122), .Y(n10117) );
  CLKINVX2TS U10702 ( .A(n7325), .Y(n10030) );
  NOR2X1TS U10703 ( .A(n12498), .B(n10774), .Y(n4099) );
  INVX1TS U10704 ( .A(n12416), .Y(n9731) );
  CLKINVX2TS U10705 ( .A(n7314), .Y(n10646) );
  CLKINVX2TS U10706 ( .A(n10814), .Y(n10861) );
  INVX1TS U10707 ( .A(n5461), .Y(n11247) );
  CLKBUFX2TS U10708 ( .A(n11591), .Y(n7339) );
  INVX2TS U10709 ( .A(n9861), .Y(n11551) );
  NOR2X1TS U10710 ( .A(n12489), .B(n12616), .Y(n7834) );
  INVX1TS U10711 ( .A(n7827), .Y(n12190) );
  INVX2TS U10712 ( .A(n4482), .Y(n10134) );
  CLKBUFX2TS U10713 ( .A(n11150), .Y(n7315) );
  INVX2TS U10714 ( .A(n3772), .Y(n11309) );
  INVX2TS U10715 ( .A(n12426), .Y(n9734) );
  INVX2TS U10716 ( .A(n7733), .Y(n10082) );
  AOI22X1TS U10717 ( .A0(n11821), .A1(n2978), .B0(n12645), .B1(n12332), .Y(
        n3101) );
  INVX1TS U10718 ( .A(n7827), .Y(n12191) );
  INVX2TS U10719 ( .A(n11144), .Y(n11107) );
  INVX1TS U10720 ( .A(n1691), .Y(n12181) );
  INVX2TS U10721 ( .A(n10388), .Y(n11727) );
  AOI211X1TS U10722 ( .A0(n10296), .A1(n12365), .B0(n2242), .C0(n2710), .Y(
        n2439) );
  AOI22X1TS U10723 ( .A0(n10070), .A1(n12489), .B0(n12634), .B1(n11096), .Y(
        n8292) );
  INVX2TS U10724 ( .A(n7733), .Y(n10081) );
  INVX1TS U10725 ( .A(n9861), .Y(n11553) );
  AOI22X1TS U10726 ( .A0(n11914), .A1(n10281), .B0(n11956), .B1(n11098), .Y(
        n8023) );
  INVX2TS U10727 ( .A(n3500), .Y(n11803) );
  CLKINVX2TS U10728 ( .A(n10477), .Y(n10810) );
  CLKINVX1TS U10729 ( .A(n11146), .Y(n11108) );
  INVX2TS U10730 ( .A(n5479), .Y(n11687) );
  INVX2TS U10731 ( .A(n12406), .Y(n9646) );
  INVX2TS U10732 ( .A(n7651), .Y(n12364) );
  INVX2TS U10733 ( .A(n3772), .Y(n11308) );
  INVX2TS U10734 ( .A(n7325), .Y(n10029) );
  INVX2TS U10735 ( .A(n8270), .Y(n9628) );
  INVX2TS U10736 ( .A(n7827), .Y(n12189) );
  INVX1TS U10737 ( .A(n11590), .Y(n10615) );
  INVX2TS U10738 ( .A(n4506), .Y(n9679) );
  INVX2TS U10739 ( .A(n9862), .Y(n11552) );
  INVX2TS U10740 ( .A(n9501), .Y(n12552) );
  INVX2TS U10741 ( .A(n10495), .Y(n10838) );
  NOR2X1TS U10742 ( .A(n12514), .B(n10762), .Y(n4043) );
  AOI22X1TS U10743 ( .A0(n12421), .A1(n10774), .B0(n11280), .B1(n12508), .Y(
        n4700) );
  INVX2TS U10744 ( .A(n10475), .Y(n10809) );
  INVX2TS U10745 ( .A(n7167), .Y(n11826) );
  INVX2TS U10746 ( .A(n7167), .Y(n11824) );
  OAI21X1TS U10747 ( .A0(n11813), .A1(n11635), .B0(n9889), .Y(n8166) );
  AOI22X1TS U10748 ( .A0(n12591), .A1(n11223), .B0(n11700), .B1(n12519), .Y(
        n5503) );
  INVX2TS U10749 ( .A(n3724), .Y(n11745) );
  INVX2TS U10750 ( .A(n12404), .Y(n9647) );
  CLKINVX2TS U10751 ( .A(n10439), .Y(n10929) );
  AOI22X1TS U10752 ( .A0(n12409), .A1(n11008), .B0(n11325), .B1(n12520), .Y(
        n6500) );
  INVX2TS U10753 ( .A(n10537), .Y(n11705) );
  INVX2TS U10754 ( .A(n1691), .Y(n12180) );
  OAI21X1TS U10755 ( .A0(n11616), .A1(n11140), .B0(n12488), .Y(n8459) );
  INVX2TS U10756 ( .A(n3706), .Y(n11356) );
  INVX2TS U10757 ( .A(n7231), .Y(n12314) );
  AOI22X1TS U10758 ( .A0(n11192), .A1(n12479), .B0(n12342), .B1(n11092), .Y(
        n8510) );
  INVX2TS U10759 ( .A(n2040), .Y(n9959) );
  INVX2TS U10760 ( .A(n12101), .Y(n11479) );
  INVX2TS U10761 ( .A(n3724), .Y(n11743) );
  INVX2TS U10762 ( .A(n7229), .Y(n10017) );
  CLKINVX2TS U10763 ( .A(n2041), .Y(n10606) );
  INVX2TS U10764 ( .A(n12103), .Y(n11480) );
  INVX2TS U10765 ( .A(n5922), .Y(n10221) );
  INVX2TS U10766 ( .A(n10389), .Y(n11726) );
  AOI22X1TS U10767 ( .A0(n11768), .A1(n10812), .B0(n12201), .B1(n11375), .Y(
        n5075) );
  INVX2TS U10768 ( .A(n5461), .Y(n11246) );
  CLKINVX2TS U10769 ( .A(n3500), .Y(n11805) );
  CLKINVX2TS U10770 ( .A(n12030), .Y(n10454) );
  INVX2TS U10771 ( .A(n10422), .Y(n10904) );
  INVX2TS U10772 ( .A(n7157), .Y(n10269) );
  AOI22X1TS U10773 ( .A0(n12342), .A1(n8211), .B0(n11504), .B1(n12134), .Y(
        n8484) );
  INVX2TS U10774 ( .A(n3724), .Y(n11744) );
  AOI22X1TS U10775 ( .A0(n11716), .A1(n5677), .B0(n11998), .B1(n11760), .Y(
        n6634) );
  INVX1TS U10776 ( .A(n3706), .Y(n11358) );
  AOI22X1TS U10777 ( .A0(n11463), .A1(n11053), .B0(n11061), .B1(n10014), .Y(
        n7183) );
  INVX2TS U10778 ( .A(n9500), .Y(n12551) );
  INVX1TS U10779 ( .A(n9500), .Y(n12550) );
  INVX2TS U10780 ( .A(n7167), .Y(n11825) );
  INVX2TS U10781 ( .A(n7157), .Y(n10270) );
  INVX2TS U10782 ( .A(n5527), .Y(n11294) );
  OAI31X1TS U10783 ( .A0(n10583), .A1(n12326), .A2(n2577), .B0(n12648), .Y(
        n2597) );
  AOI22X1TS U10784 ( .A0(n11839), .A1(n2122), .B0(n9725), .B1(n2124), .Y(n2117) );
  INVX2TS U10785 ( .A(n5527), .Y(n11293) );
  AOI22X1TS U10786 ( .A0(n5770), .A1(n10577), .B0(n11348), .B1(n11759), .Y(
        n6642) );
  INVX1TS U10787 ( .A(n5527), .Y(n11295) );
  OAI31X1TS U10788 ( .A0(n12345), .A1(n11491), .A2(n12135), .B0(n11946), .Y(
        n7959) );
  CLKINVX2TS U10789 ( .A(n7293), .Y(n9487) );
  AOI22X1TS U10790 ( .A0(n12288), .A1(n12614), .B0(n10589), .B1(n11068), .Y(
        n2625) );
  INVX2TS U10791 ( .A(n5922), .Y(n10222) );
  INVX2TS U10792 ( .A(n12424), .Y(n9735) );
  AOI22X1TS U10793 ( .A0(n11579), .A1(n12343), .B0(n11192), .B1(n9481), .Y(
        n8253) );
  INVX2TS U10794 ( .A(n10536), .Y(n11706) );
  INVX2TS U10795 ( .A(n7293), .Y(n9486) );
  AOI22X1TS U10796 ( .A0(n12343), .A1(n10643), .B0(n12478), .B1(n12471), .Y(
        n8496) );
  INVX1TS U10797 ( .A(n7629), .Y(n10702) );
  OR2X2TS U10798 ( .A(n12338), .B(n12289), .Y(n1956) );
  INVX2TS U10799 ( .A(n10441), .Y(n10930) );
  INVX2TS U10800 ( .A(n7629), .Y(n10701) );
  NOR2X1TS U10801 ( .A(n12526), .B(n11008), .Y(n5899) );
  INVX2TS U10802 ( .A(n8209), .Y(n10102) );
  INVX2TS U10803 ( .A(n8209), .Y(n10101) );
  CLKINVX2TS U10804 ( .A(n7276), .Y(n12129) );
  INVX2TS U10805 ( .A(n7975), .Y(n9629) );
  OAI21X1TS U10806 ( .A0(n10875), .A1(n10411), .B0(n12017), .Y(n4813) );
  OAI21X1TS U10807 ( .A0(n10798), .A1(n10415), .B0(n11781), .Y(n4812) );
  INVX2TS U10808 ( .A(n4066), .Y(n10109) );
  AOI22X1TS U10809 ( .A0(n11789), .A1(n11814), .B0(n11027), .B1(n10013), .Y(
        n8626) );
  INVX2TS U10810 ( .A(n7893), .Y(n11160) );
  AOI22X1TS U10811 ( .A0(n2611), .A1(n11422), .B0(n11918), .B1(n11518), .Y(
        n2985) );
  INVX2TS U10812 ( .A(n10535), .Y(n11704) );
  INVX2TS U10813 ( .A(n7893), .Y(n11159) );
  INVX2TS U10814 ( .A(n4575), .Y(n9691) );
  INVX1TS U10815 ( .A(n12100), .Y(n11481) );
  INVX2TS U10816 ( .A(n3706), .Y(n11357) );
  AOI22X1TS U10817 ( .A0(n11769), .A1(n11781), .B0(n11701), .B1(n12029), .Y(
        n4871) );
  INVX1TS U10818 ( .A(n7231), .Y(n12312) );
  AOI22X1TS U10819 ( .A0(n11249), .A1(n10401), .B0(n11779), .B1(n10411), .Y(
        n4562) );
  CLKINVX2TS U10820 ( .A(n2040), .Y(n9960) );
  INVX2TS U10821 ( .A(n11588), .Y(n10616) );
  AOI22X1TS U10822 ( .A0(n11821), .A1(n10171), .B0(n12324), .B1(n11514), .Y(
        n2553) );
  INVX1TS U10823 ( .A(n1691), .Y(n12182) );
  OAI31X1TS U10824 ( .A0(n11716), .A1(n12280), .A2(n11999), .B0(n11722), .Y(
        n5592) );
  AOI22X1TS U10825 ( .A0(n11506), .A1(n2518), .B0(n11453), .B1(n2185), .Y(
        n2543) );
  AOI22X1TS U10826 ( .A0(n11767), .A1(n12029), .B0(n11375), .B1(n12016), .Y(
        n5086) );
  AOI22X1TS U10827 ( .A0(n12437), .A1(n10762), .B0(n11328), .B1(n12523), .Y(
        n4628) );
  CLKINVX2TS U10828 ( .A(n10813), .Y(n10860) );
  CLKINVX2TS U10829 ( .A(n10423), .Y(n10903) );
  INVX2TS U10830 ( .A(n12418), .Y(n9730) );
  INVX2TS U10831 ( .A(n5479), .Y(n11686) );
  CLKINVX2TS U10832 ( .A(n3518), .Y(n10922) );
  INVX2TS U10833 ( .A(n4482), .Y(n10133) );
  NOR2X1TS U10834 ( .A(n12510), .B(n10996), .Y(n5843) );
  INVX1TS U10835 ( .A(n3772), .Y(n11310) );
  INVX2TS U10836 ( .A(n5479), .Y(n11688) );
  AOI22X1TS U10837 ( .A0(n12393), .A1(n10996), .B0(n11277), .B1(n12504), .Y(
        n6428) );
  CLKINVX2TS U10838 ( .A(n5316), .Y(n10847) );
  CLKINVX2TS U10839 ( .A(n4066), .Y(n10110) );
  CLKINVX2TS U10840 ( .A(n5298), .Y(n11691) );
  INVX2TS U10841 ( .A(n4575), .Y(n9690) );
  INVX2TS U10842 ( .A(n4506), .Y(n9680) );
  OAI31X1TS U10843 ( .A0(n12217), .A1(n12233), .A2(n10457), .B0(n12226), .Y(
        n5439) );
  INVX2TS U10844 ( .A(n4122), .Y(n10118) );
  INVX2TS U10845 ( .A(n5866), .Y(n10214) );
  INVX2TS U10846 ( .A(n5866), .Y(n10213) );
  AOI22X1TS U10847 ( .A0(n12582), .A1(n11211), .B0(n11682), .B1(n12502), .Y(
        n5437) );
  INVX2TS U10848 ( .A(n5461), .Y(n11245) );
  CLKINVX2TS U10849 ( .A(n10493), .Y(n10837) );
  INVX2TS U10850 ( .A(n5316), .Y(n10846) );
  CLKINVX2TS U10851 ( .A(n3500), .Y(n11804) );
  CLKINVX2TS U10852 ( .A(n5298), .Y(n11690) );
  INVX2TS U10853 ( .A(n9501), .Y(n12553) );
  INVX2TS U10854 ( .A(n5600), .Y(n10488) );
  CLKINVX2TS U10855 ( .A(n10813), .Y(n10859) );
  CLKBUFX2TS U10856 ( .A(n11746), .Y(n5658) );
  CLKINVX2TS U10857 ( .A(n5750), .Y(n11747) );
  INVX1TS U10858 ( .A(n9402), .Y(n11997) );
  INVX1TS U10859 ( .A(n10529), .Y(n12224) );
  CLKINVX2TS U10860 ( .A(n4130), .Y(n9147) );
  INVX2TS U10861 ( .A(n3761), .Y(n9110) );
  INVX2TS U10862 ( .A(n10711), .Y(n10282) );
  INVX1TS U10863 ( .A(n7310), .Y(n11097) );
  INVX2TS U10864 ( .A(n9809), .Y(n11788) );
  INVX2TS U10865 ( .A(n5577), .Y(n12431) );
  CLKINVX2TS U10866 ( .A(n2358), .Y(n12080) );
  INVX2TS U10867 ( .A(n5900), .Y(n11389) );
  CLKINVX2TS U10868 ( .A(n11277), .Y(n10428) );
  INVX1TS U10869 ( .A(n7815), .Y(n10729) );
  INVX2TS U10870 ( .A(n8231), .Y(n11192) );
  INVX2TS U10871 ( .A(n11993), .Y(n11732) );
  INVX2TS U10872 ( .A(n1811), .Y(n11917) );
  INVX1TS U10873 ( .A(n6320), .Y(n10576) );
  NOR2X1TS U10874 ( .A(n10585), .B(n12408), .Y(n5719) );
  CLKINVX2TS U10875 ( .A(n5761), .Y(n11371) );
  CLKINVX2TS U10876 ( .A(n1875), .Y(n12352) );
  INVX2TS U10877 ( .A(n11423), .Y(n10007) );
  CLKBUFX2TS U10878 ( .A(n10966), .Y(n1986) );
  INVX2TS U10879 ( .A(n11994), .Y(n11733) );
  CLKINVX2TS U10880 ( .A(n2061), .Y(n12118) );
  INVX2TS U10881 ( .A(n3662), .Y(n11768) );
  INVX2TS U10882 ( .A(n5514), .Y(n11699) );
  CLKBUFX2TS U10883 ( .A(n9923), .Y(n1968) );
  INVX2TS U10884 ( .A(n3579), .Y(n10887) );
  INVX2TS U10885 ( .A(n12025), .Y(n11681) );
  INVX2TS U10886 ( .A(n8231), .Y(n11193) );
  INVX2TS U10887 ( .A(n10381), .Y(n12237) );
  INVX2TS U10888 ( .A(n10855), .Y(n10105) );
  INVX1TS U10889 ( .A(n12140), .Y(n12174) );
  INVX2TS U10890 ( .A(n6320), .Y(n10577) );
  INVX2TS U10891 ( .A(n6025), .Y(n9994) );
  CLKINVX2TS U10892 ( .A(n3827), .Y(n12390) );
  CLKINVX2TS U10893 ( .A(n5782), .Y(n10980) );
  INVX2TS U10894 ( .A(n2629), .Y(n12291) );
  INVX2TS U10895 ( .A(n7286), .Y(n9481) );
  INVX2TS U10896 ( .A(n10835), .Y(n10185) );
  CLKINVX2TS U10897 ( .A(n1714), .Y(n12474) );
  INVX2TS U10898 ( .A(n2252), .Y(n9079) );
  INVX1TS U10899 ( .A(n3950), .Y(n10410) );
  INVX2TS U10900 ( .A(n1811), .Y(n11919) );
  CLKINVX1TS U10901 ( .A(n1714), .Y(n12477) );
  CLKINVX1TS U10902 ( .A(n1875), .Y(n12354) );
  INVX2TS U10903 ( .A(n5338), .Y(n10863) );
  INVX1TS U10904 ( .A(n12232), .Y(n10505) );
  AOI22X1TS U10905 ( .A0(n12245), .A1(n11393), .B0(n10899), .B1(n12501), .Y(
        n4189) );
  INVX2TS U10906 ( .A(n5377), .Y(n10880) );
  CLKINVX2TS U10907 ( .A(n3695), .Y(n9103) );
  INVX2TS U10908 ( .A(n2413), .Y(n10203) );
  INVX2TS U10909 ( .A(n2171), .Y(n11524) );
  CLKINVX2TS U10910 ( .A(n5622), .Y(n12441) );
  INVX2TS U10911 ( .A(n10885), .Y(n10209) );
  INVX2TS U10912 ( .A(n1712), .Y(n11625) );
  INVX1TS U10913 ( .A(n10631), .Y(n10949) );
  INVX2TS U10914 ( .A(n10531), .Y(n12225) );
  INVX2TS U10915 ( .A(n5338), .Y(n10862) );
  NOR2X1TS U10916 ( .A(n12235), .B(n11000), .Y(n6433) );
  INVX1TS U10917 ( .A(n10383), .Y(n12238) );
  INVX2TS U10918 ( .A(n3926), .Y(n10414) );
  INVX2TS U10919 ( .A(n10885), .Y(n10210) );
  INVX1TS U10920 ( .A(n7233), .Y(n11475) );
  INVX2TS U10921 ( .A(n9677), .Y(n11212) );
  INVX1TS U10922 ( .A(n12380), .Y(n9175) );
  INVX2TS U10923 ( .A(n1886), .Y(n9112) );
  INVX2TS U10924 ( .A(n10867), .Y(n10806) );
  INVX2TS U10925 ( .A(n3693), .Y(n11751) );
  CLKBUFX2TS U10926 ( .A(n3930), .Y(n12566) );
  INVX1TS U10927 ( .A(n3644), .Y(n10877) );
  INVX2TS U10928 ( .A(n1752), .Y(n12458) );
  INVX1TS U10929 ( .A(n10529), .Y(n12227) );
  NOR2X1TS U10930 ( .A(n10408), .B(n12420), .Y(n3889) );
  CLKINVX1TS U10931 ( .A(n1712), .Y(n11626) );
  INVX2TS U10932 ( .A(n11102), .Y(n11915) );
  CLKINVX2TS U10933 ( .A(n12138), .Y(n12175) );
  INVX2TS U10934 ( .A(n3930), .Y(n12569) );
  INVX2TS U10935 ( .A(n10541), .Y(n12248) );
  INVX2TS U10936 ( .A(n9673), .Y(n11702) );
  INVX1TS U10937 ( .A(n10540), .Y(n12250) );
  INVX2TS U10938 ( .A(n3531), .Y(n10489) );
  INVX2TS U10939 ( .A(n12120), .Y(n10321) );
  INVX2TS U10940 ( .A(n3662), .Y(n11767) );
  CLKINVX2TS U10941 ( .A(n11003), .Y(n9995) );
  NOR2X1TS U10942 ( .A(n12419), .B(n11321), .Y(n4459) );
  INVX2TS U10943 ( .A(n7815), .Y(n10728) );
  INVX2TS U10944 ( .A(n12154), .Y(n9968) );
  INVX2TS U10945 ( .A(n1750), .Y(n11607) );
  INVX2TS U10946 ( .A(n9781), .Y(n11349) );
  INVX1TS U10947 ( .A(n7666), .Y(n11593) );
  INVX1TS U10948 ( .A(n5377), .Y(n10879) );
  CLKINVX2TS U10949 ( .A(n12235), .Y(n10506) );
  INVX2TS U10950 ( .A(n12068), .Y(n9576) );
  CLKINVX2TS U10951 ( .A(n12254), .Y(n10425) );
  OAI31X1TS U10952 ( .A0(n11911), .A1(n12358), .A2(n11595), .B0(n12647), .Y(
        n2582) );
  CLKINVX2TS U10953 ( .A(n2358), .Y(n12078) );
  INVX1TS U10954 ( .A(n7476), .Y(n12618) );
  INVX2TS U10955 ( .A(n2629), .Y(n12288) );
  OAI21X1TS U10956 ( .A0(n11022), .A1(n12652), .B0(n10223), .Y(n3048) );
  CLKINVX2TS U10957 ( .A(n1711), .Y(n12483) );
  INVX2TS U10958 ( .A(n12068), .Y(n9575) );
  INVX1TS U10959 ( .A(n8231), .Y(n11194) );
  INVX1TS U10960 ( .A(n7185), .Y(n11055) );
  CLKINVX2TS U10961 ( .A(n1750), .Y(n11606) );
  INVX1TS U10962 ( .A(n9552), .Y(n12350) );
  INVX2TS U10963 ( .A(n3912), .Y(n11250) );
  INVX1TS U10964 ( .A(n12209), .Y(n9970) );
  INVX2TS U10965 ( .A(n2562), .Y(n10172) );
  INVX2TS U10966 ( .A(n2319), .Y(n9072) );
  INVX1TS U10967 ( .A(n5506), .Y(n10466) );
  CLKINVX2TS U10968 ( .A(n9091), .Y(n12116) );
  INVX1TS U10969 ( .A(n9701), .Y(n11158) );
  NOR2X1TS U10970 ( .A(n12254), .B(n10766), .Y(n4633) );
  INVX2TS U10971 ( .A(n7390), .Y(n10668) );
  INVX1TS U10972 ( .A(n7390), .Y(n10670) );
  CLKINVX2TS U10973 ( .A(n11596), .Y(n9964) );
  AOI22X1TS U10974 ( .A0(n12241), .A1(n11222), .B0(n10868), .B1(n12529), .Y(
        n6099) );
  INVX2TS U10975 ( .A(n3579), .Y(n10888) );
  INVX2TS U10976 ( .A(n12138), .Y(n12173) );
  CLKINVX1TS U10977 ( .A(n4296), .Y(n10790) );
  INVX1TS U10978 ( .A(n10394), .Y(n12261) );
  INVX2TS U10979 ( .A(n3644), .Y(n10876) );
  INVX2TS U10980 ( .A(n7185), .Y(n11053) );
  CLKINVX2TS U10981 ( .A(n5900), .Y(n11390) );
  INVX2TS U10982 ( .A(n3671), .Y(n12022) );
  CLKINVX2TS U10983 ( .A(n11031), .Y(n11070) );
  INVX2TS U10984 ( .A(n5844), .Y(n11384) );
  INVX2TS U10985 ( .A(n11611), .Y(n9870) );
  CLKINVX2TS U10986 ( .A(n1755), .Y(n11127) );
  INVX2TS U10987 ( .A(n3540), .Y(n10905) );
  CLKINVX2TS U10988 ( .A(n10514), .Y(n11015) );
  INVX2TS U10989 ( .A(n1712), .Y(n11624) );
  INVX1TS U10990 ( .A(n5440), .Y(n10458) );
  INVX2TS U10991 ( .A(n7692), .Y(n9543) );
  INVX1TS U10992 ( .A(n10042), .Y(n11066) );
  CLKINVX2TS U10993 ( .A(n2171), .Y(n11526) );
  AOI22X1TS U10994 ( .A0(n12218), .A1(n11210), .B0(n10851), .B1(n12513), .Y(
        n6055) );
  INVX1TS U10995 ( .A(n7725), .Y(n11151) );
  CLKINVX2TS U10996 ( .A(n3761), .Y(n9111) );
  INVX2TS U10997 ( .A(n7724), .Y(n9866) );
  AOI22X1TS U10998 ( .A0(n10169), .A1(n11014), .B0(n12528), .B1(n11283), .Y(
        n6817) );
  INVX2TS U10999 ( .A(n10933), .Y(n10123) );
  CLKINVX2TS U11000 ( .A(n1711), .Y(n12484) );
  CLKINVX2TS U11001 ( .A(n12311), .Y(n11036) );
  CLKINVX1TS U11002 ( .A(n4013), .Y(n10758) );
  INVX2TS U11003 ( .A(n4119), .Y(n10114) );
  CLKINVX2TS U11004 ( .A(n5953), .Y(n11018) );
  CLKINVX2TS U11005 ( .A(n2061), .Y(n12117) );
  INVX2TS U11006 ( .A(n8159), .Y(n9890) );
  INVX2TS U11007 ( .A(n11521), .Y(n10069) );
  INVX2TS U11008 ( .A(n4100), .Y(n11236) );
  CLKINVX2TS U11009 ( .A(n11068), .Y(n10593) );
  CLKINVX2TS U11010 ( .A(n3827), .Y(n12389) );
  INVX1TS U11011 ( .A(n4013), .Y(n10759) );
  CLKINVX2TS U11012 ( .A(n12310), .Y(n11034) );
  CLKINVX2TS U11013 ( .A(n5450), .Y(n9293) );
  INVX2TS U11014 ( .A(n3662), .Y(n11769) );
  INVX2TS U11015 ( .A(n7281), .Y(n10639) );
  INVX2TS U11016 ( .A(n10924), .Y(n11008) );
  INVX2TS U11017 ( .A(n3490), .Y(n11809) );
  AOI22X1TS U11018 ( .A0(n10161), .A1(n11002), .B0(n12513), .B1(n11233), .Y(
        n6759) );
  CLKINVX2TS U11019 ( .A(n3630), .Y(n12038) );
  INVX2TS U11020 ( .A(n3950), .Y(n10411) );
  INVX2TS U11021 ( .A(n12120), .Y(n10320) );
  INVX2TS U11022 ( .A(n7473), .Y(n11898) );
  INVX1TS U11023 ( .A(n5338), .Y(n10864) );
  INVX2TS U11024 ( .A(n5577), .Y(n12432) );
  INVX2TS U11025 ( .A(n3490), .Y(n11811) );
  INVX2TS U11026 ( .A(n10896), .Y(n10995) );
  CLKINVX2TS U11027 ( .A(n10613), .Y(n10664) );
  INVX2TS U11028 ( .A(n10866), .Y(n10808) );
  INVX2TS U11029 ( .A(n10897), .Y(n10996) );
  INVX2TS U11030 ( .A(n12375), .Y(n10119) );
  INVX2TS U11031 ( .A(n3827), .Y(n12387) );
  INVX2TS U11032 ( .A(n9782), .Y(n11348) );
  NOR2X1TS U11033 ( .A(n12409), .B(n11282), .Y(n6262) );
  INVX2TS U11034 ( .A(n3498), .Y(n9919) );
  INVX2TS U11035 ( .A(n11386), .Y(n10121) );
  INVX2TS U11036 ( .A(n3486), .Y(n10163) );
  CLKINVX2TS U11037 ( .A(n4044), .Y(n11244) );
  INVX2TS U11038 ( .A(n10629), .Y(n10948) );
  INVX2TS U11039 ( .A(n4013), .Y(n10757) );
  CLKINVX2TS U11040 ( .A(n5750), .Y(n11748) );
  CLKINVX2TS U11041 ( .A(n1752), .Y(n12460) );
  CLKINVX2TS U11042 ( .A(n7066), .Y(n9463) );
  INVX1TS U11043 ( .A(n11535), .Y(n9838) );
  INVX2TS U11044 ( .A(n2413), .Y(n10204) );
  INVX2TS U11045 ( .A(n5671), .Y(n11354) );
  INVX2TS U11046 ( .A(n3926), .Y(n10415) );
  INVX1TS U11047 ( .A(n5671), .Y(n11355) );
  INVX2TS U11048 ( .A(n9403), .Y(n11998) );
  CLKINVX2TS U11049 ( .A(n12378), .Y(n10120) );
  INVX2TS U11050 ( .A(n2145), .Y(n11827) );
  INVX2TS U11051 ( .A(n5953), .Y(n11019) );
  CLKINVX2TS U11052 ( .A(n3498), .Y(n9920) );
  INVX2TS U11053 ( .A(n3841), .Y(n9917) );
  INVX2TS U11054 ( .A(n10923), .Y(n11007) );
  INVX2TS U11055 ( .A(n12145), .Y(n10207) );
  INVX2TS U11056 ( .A(n10630), .Y(n10950) );
  INVX2TS U11057 ( .A(n11990), .Y(n10202) );
  CLKINVX2TS U11058 ( .A(n1974), .Y(n11074) );
  INVX2TS U11059 ( .A(n12447), .Y(n10189) );
  CLKINVX1TS U11060 ( .A(n1886), .Y(n9113) );
  CLKINVX2TS U11061 ( .A(n5516), .Y(n9303) );
  INVX1TS U11062 ( .A(n5577), .Y(n12434) );
  INVX2TS U11063 ( .A(n7458), .Y(n10302) );
  INVX1TS U11064 ( .A(n5440), .Y(n10457) );
  AOI22X1TS U11065 ( .A0(n11341), .A1(n11981), .B0(n11697), .B1(n12574), .Y(
        n6556) );
  INVX2TS U11066 ( .A(n12626), .Y(n10347) );
  AOI22X1TS U11067 ( .A0(n12340), .A1(n10227), .B0(n11040), .B1(n12454), .Y(
        n3062) );
  INVX2TS U11068 ( .A(n9678), .Y(n11214) );
  INVX2TS U11069 ( .A(n2312), .Y(n10977) );
  INVX2TS U11070 ( .A(n7692), .Y(n9542) );
  CLKINVX2TS U11071 ( .A(n5874), .Y(n9330) );
  CLKINVX2TS U11072 ( .A(n10831), .Y(n9135) );
  CLKINVX2TS U11073 ( .A(n1711), .Y(n12485) );
  INVX2TS U11074 ( .A(n5750), .Y(n11746) );
  CLKINVX2TS U11075 ( .A(n10935), .Y(n9346) );
  INVX2TS U11076 ( .A(n7693), .Y(n11139) );
  INVX2TS U11077 ( .A(n5622), .Y(n12439) );
  INVX2TS U11078 ( .A(n5296), .Y(n9941) );
  AOI22X1TS U11079 ( .A0(n10967), .A1(n10196), .B0(n12112), .B1(n12453), .Y(
        n3063) );
  INVX2TS U11080 ( .A(n6025), .Y(n9993) );
  CLKINVX2TS U11081 ( .A(n2312), .Y(n10978) );
  NOR2X1TS U11082 ( .A(n12394), .B(n11234), .Y(n6222) );
  INVX2TS U11083 ( .A(n3644), .Y(n10875) );
  CLKINVX1TS U11084 ( .A(n4100), .Y(n11238) );
  CLKINVX1TS U11085 ( .A(n3930), .Y(n12567) );
  CLKINVX2TS U11086 ( .A(n11325), .Y(n10445) );
  INVX2TS U11087 ( .A(n5798), .Y(n10983) );
  INVX2TS U11088 ( .A(n7476), .Y(n12617) );
  CLKINVX2TS U11089 ( .A(n12253), .Y(n10426) );
  INVX2TS U11090 ( .A(n9673), .Y(n11701) );
  INVX2TS U11091 ( .A(n5844), .Y(n11383) );
  NOR2X1TS U11092 ( .A(n12231), .B(n10779), .Y(n4705) );
  INVX2TS U11093 ( .A(n5761), .Y(n11372) );
  INVX1TS U11094 ( .A(n3693), .Y(n11749) );
  INVX2TS U11095 ( .A(n2457), .Y(n10199) );
  INVX2TS U11096 ( .A(n5577), .Y(n12433) );
  CLKINVX2TS U11097 ( .A(n1702), .Y(n10676) );
  INVX2TS U11098 ( .A(n2145), .Y(n11829) );
  INVX2TS U11099 ( .A(n12344), .Y(n11586) );
  INVX2TS U11100 ( .A(n3540), .Y(n10907) );
  INVX2TS U11101 ( .A(n1875), .Y(n12353) );
  INVX2TS U11102 ( .A(n9677), .Y(n11213) );
  INVX2TS U11103 ( .A(n7473), .Y(n11897) );
  INVX2TS U11104 ( .A(n7476), .Y(n12616) );
  CLKINVX2TS U11105 ( .A(n1711), .Y(n12482) );
  INVX2TS U11106 ( .A(n2629), .Y(n12289) );
  CLKINVX2TS U11107 ( .A(n8191), .Y(n11183) );
  INVX2TS U11108 ( .A(n12212), .Y(n9969) );
  INVX2TS U11109 ( .A(n5450), .Y(n9292) );
  INVX2TS U11110 ( .A(n12626), .Y(n10346) );
  INVX2TS U11111 ( .A(n11609), .Y(n9869) );
  INVX1TS U11112 ( .A(n7473), .Y(n11896) );
  INVX2TS U11113 ( .A(n9552), .Y(n12351) );
  INVX1TS U11114 ( .A(n10530), .Y(n12226) );
  INVX2TS U11115 ( .A(n11388), .Y(n10122) );
  INVX1TS U11116 ( .A(n11177), .Y(n11497) );
  INVX2TS U11117 ( .A(n12234), .Y(n10507) );
  INVX2TS U11118 ( .A(n10094), .Y(n11133) );
  CLKINVX2TS U11119 ( .A(n11067), .Y(n10592) );
  NOR2X1TS U11120 ( .A(n10581), .B(n12392), .Y(n5694) );
  CLKINVX2TS U11121 ( .A(n10532), .Y(n11147) );
  INVX2TS U11122 ( .A(n12228), .Y(n10418) );
  INVX2TS U11123 ( .A(n7233), .Y(n11474) );
  INVX2TS U11124 ( .A(n10711), .Y(n10281) );
  INVX2TS U11125 ( .A(n11178), .Y(n11499) );
  INVX2TS U11126 ( .A(n5514), .Y(n11700) );
  CLKINVX2TS U11127 ( .A(n10516), .Y(n11016) );
  INVX1TS U11128 ( .A(n12255), .Y(n10511) );
  INVX1TS U11129 ( .A(n10392), .Y(n12259) );
  CLKINVX2TS U11130 ( .A(n4044), .Y(n11243) );
  INVX2TS U11131 ( .A(n3912), .Y(n11249) );
  INVX1TS U11132 ( .A(n10542), .Y(n12249) );
  AOI22X1TS U11133 ( .A0(n10135), .A1(n10768), .B0(n12516), .B1(n11370), .Y(
        n4960) );
  INVX2TS U11134 ( .A(n8159), .Y(n9889) );
  CLKINVX1TS U11135 ( .A(n1749), .Y(n12469) );
  CLKINVX2TS U11136 ( .A(n2291), .Y(n12087) );
  INVX2TS U11137 ( .A(n11594), .Y(n9963) );
  INVX2TS U11138 ( .A(n10381), .Y(n12236) );
  CLKINVX2TS U11139 ( .A(n5622), .Y(n12442) );
  CLKINVX2TS U11140 ( .A(n1752), .Y(n12459) );
  INVX2TS U11141 ( .A(n4119), .Y(n10113) );
  AOI22X1TS U11142 ( .A0(n12268), .A1(n11405), .B0(n10915), .B1(n12517), .Y(
        n4145) );
  CLKINVX2TS U11143 ( .A(n11029), .Y(n11853) );
  INVX2TS U11144 ( .A(n5516), .Y(n9302) );
  CLKINVX2TS U11145 ( .A(n1755), .Y(n11126) );
  INVX2TS U11146 ( .A(n2245), .Y(n10992) );
  INVX1TS U11147 ( .A(n10382), .Y(n12239) );
  INVX2TS U11148 ( .A(n8093), .Y(n9885) );
  AOI32XLTS U11149 ( .A0(n3830), .A1(n12046), .A2(sa33[4]), .B0(n10126), .B1(
        n12044), .Y(n4357) );
  INVX2TS U11150 ( .A(n10843), .Y(n10761) );
  INVX2TS U11151 ( .A(n9810), .Y(n11789) );
  INVX2TS U11152 ( .A(n9674), .Y(n11703) );
  INVX2TS U11153 ( .A(n7725), .Y(n11150) );
  INVX1TS U11154 ( .A(n3841), .Y(n9918) );
  INVX1TS U11155 ( .A(n7390), .Y(n10669) );
  INVX2TS U11156 ( .A(n10845), .Y(n10762) );
  INVX2TS U11157 ( .A(n7458), .Y(n10301) );
  INVX2TS U11158 ( .A(n2457), .Y(n10200) );
  AOI22X1TS U11159 ( .A0(n11042), .A1(n11068), .B0(n12652), .B1(n10196), .Y(
        n2754) );
  INVX2TS U11160 ( .A(n12132), .Y(n10216) );
  INVX1TS U11161 ( .A(n3579), .Y(n10889) );
  INVX2TS U11162 ( .A(n12163), .Y(n10089) );
  INVX2TS U11163 ( .A(n10041), .Y(n11065) );
  INVX1TS U11164 ( .A(n7693), .Y(n11140) );
  CLKINVX2TS U11165 ( .A(n12125), .Y(n12166) );
  INVX2TS U11166 ( .A(n10865), .Y(n10807) );
  INVX1TS U11167 ( .A(n7281), .Y(n10638) );
  INVX2TS U11168 ( .A(n7299), .Y(n12481) );
  INVX1TS U11169 ( .A(n7292), .Y(n12135) );
  CLKINVX2TS U11170 ( .A(n1740), .Y(n10663) );
  INVX2TS U11171 ( .A(n7737), .Y(n11156) );
  INVX1TS U11172 ( .A(n7666), .Y(n11592) );
  INVX2TS U11173 ( .A(n5671), .Y(n11353) );
  INVX2TS U11174 ( .A(n7299), .Y(n12478) );
  OAI21X1TS U11175 ( .A0(n10841), .A1(n12574), .B0(n10241), .Y(n6037) );
  INVX1TS U11176 ( .A(n11647), .Y(n10692) );
  CLKINVX1TS U11177 ( .A(n12231), .Y(n10419) );
  CLKINVX2TS U11178 ( .A(n12151), .Y(n9967) );
  INVX2TS U11179 ( .A(n3912), .Y(n11248) );
  AOI22X1TS U11180 ( .A0(n10128), .A1(n10779), .B0(n12499), .B1(n11321), .Y(
        n5018) );
  CLKINVX2TS U11181 ( .A(n5900), .Y(n11391) );
  INVX1TS U11182 ( .A(n10392), .Y(n12262) );
  CLKBUFX2TS U11183 ( .A(n12160), .Y(n1689) );
  INVX2TS U11184 ( .A(n12230), .Y(n10420) );
  CLKINVX2TS U11185 ( .A(n11056), .Y(n11947) );
  INVX2TS U11186 ( .A(n11101), .Y(n11914) );
  INVX2TS U11187 ( .A(n10913), .Y(n10218) );
  INVX2TS U11188 ( .A(n7666), .Y(n11591) );
  INVX1TS U11189 ( .A(n12335), .Y(n10633) );
  NOR2X1TS U11190 ( .A(n12258), .B(n11012), .Y(n6505) );
  INVX2TS U11191 ( .A(n4044), .Y(n11242) );
  INVX2TS U11192 ( .A(n7233), .Y(n11473) );
  NOR2X1TS U11193 ( .A(n10374), .B(n9634), .Y(n3507) );
  INVX2TS U11194 ( .A(n8093), .Y(n9886) );
  CLKINVX2TS U11195 ( .A(n12125), .Y(n12168) );
  NOR2X1TS U11196 ( .A(n12437), .B(n11369), .Y(n4419) );
  INVX2TS U11197 ( .A(n7737), .Y(n11155) );
  INVX2TS U11198 ( .A(n3685), .Y(n10450) );
  CLKINVX2TS U11199 ( .A(n12124), .Y(n12169) );
  INVX2TS U11200 ( .A(n11005), .Y(n9996) );
  INVX2TS U11201 ( .A(n9782), .Y(n11347) );
  CLKINVX1TS U11202 ( .A(n3671), .Y(n12023) );
  INVX2TS U11203 ( .A(n11523), .Y(n10070) );
  CLKINVX2TS U11204 ( .A(n1749), .Y(n12466) );
  INVX2TS U11205 ( .A(n3695), .Y(n9102) );
  INVX2TS U11206 ( .A(n11645), .Y(n10691) );
  INVX2TS U11207 ( .A(n2562), .Y(n10171) );
  INVX2TS U11208 ( .A(n3630), .Y(n12037) );
  AOI22X1TS U11209 ( .A0(n12648), .A1(n11004), .B0(n12154), .B1(n12091), .Y(
        n1665) );
  INVX2TS U11210 ( .A(n7310), .Y(n11096) );
  INVX2TS U11211 ( .A(n10815), .Y(n10773) );
  INVX2TS U11212 ( .A(n7292), .Y(n12136) );
  INVX2TS U11213 ( .A(n10913), .Y(n10217) );
  INVX2TS U11214 ( .A(n12337), .Y(n10632) );
  INVX2TS U11215 ( .A(n9700), .Y(n11157) );
  INVX2TS U11216 ( .A(n4100), .Y(n11237) );
  CLKINVX2TS U11217 ( .A(n1714), .Y(n12476) );
  CLKBUFX2TS U11218 ( .A(n10004), .Y(n1668) );
  INVX1TS U11219 ( .A(n3685), .Y(n10451) );
  INVX1TS U11220 ( .A(n7310), .Y(n11098) );
  INVX1TS U11221 ( .A(n12336), .Y(n10634) );
  INVX2TS U11222 ( .A(n10393), .Y(n12260) );
  INVX1TS U11223 ( .A(n5377), .Y(n10878) );
  INVX2TS U11224 ( .A(n11424), .Y(n10008) );
  INVX2TS U11225 ( .A(n8191), .Y(n11182) );
  INVX2TS U11226 ( .A(n11533), .Y(n9837) );
  INVX1TS U11227 ( .A(n10894), .Y(n10442) );
  INVX2TS U11228 ( .A(n7724), .Y(n9865) );
  CLKINVX1TS U11229 ( .A(n12126), .Y(n12167) );
  CLKINVX2TS U11230 ( .A(n1740), .Y(n10662) );
  CLKBUFX2TS U11231 ( .A(n10175), .Y(n2033) );
  NOR2X1TS U11232 ( .A(n10404), .B(n12436), .Y(n3864) );
  CLKINVX2TS U11233 ( .A(n1749), .Y(n12468) );
  OAI21X1TS U11234 ( .A0(n10927), .A1(n12592), .B0(n10125), .Y(n4270) );
  CLKINVX2TS U11235 ( .A(n1938), .Y(n12346) );
  CLKINVX1TS U11236 ( .A(n1949), .Y(n9109) );
  INVX2TS U11237 ( .A(n11176), .Y(n11498) );
  AOI22X1TS U11238 ( .A0(n11939), .A1(n11462), .B0(n11622), .B1(n7429), .Y(
        n8133) );
  INVX2TS U11239 ( .A(n1949), .Y(n9108) );
  INVX2TS U11240 ( .A(n7292), .Y(n12134) );
  INVX1TS U11241 ( .A(n3540), .Y(n10906) );
  INVX2TS U11242 ( .A(n12132), .Y(n10215) );
  INVX2TS U11243 ( .A(n7286), .Y(n9482) );
  AOI22X1TS U11244 ( .A0(n11040), .A1(n10196), .B0(n11441), .B1(n12650), .Y(
        n2647) );
  INVX2TS U11245 ( .A(n12257), .Y(n10512) );
  CLKINVX2TS U11246 ( .A(n12342), .Y(n11585) );
  INVX2TS U11247 ( .A(n4296), .Y(n10791) );
  CLKINVX2TS U11248 ( .A(n2171), .Y(n11525) );
  AOI22X1TS U11249 ( .A0(n12279), .A1(n5576), .B0(n9974), .B1(n12293), .Y(
        n5964) );
  INVX1TS U11250 ( .A(n7422), .Y(n10674) );
  INVX1TS U11251 ( .A(n9551), .Y(n12349) );
  INVX2TS U11252 ( .A(n3693), .Y(n11750) );
  INVX1TS U11253 ( .A(n10540), .Y(n12247) );
  INVX1TS U11254 ( .A(n7299), .Y(n12479) );
  AOI22X1TS U11255 ( .A0(n12370), .A1(n7665), .B0(n11958), .B1(n11124), .Y(
        n8000) );
  INVX2TS U11256 ( .A(n7422), .Y(n10673) );
  CLKINVX1TS U11257 ( .A(n1752), .Y(n12461) );
  INVX2TS U11258 ( .A(n12382), .Y(n9176) );
  INVX2TS U11259 ( .A(n7185), .Y(n11054) );
  INVX2TS U11260 ( .A(n7693), .Y(n11138) );
  INVX2TS U11261 ( .A(n12005), .Y(n10182) );
  NOR2X1TS U11262 ( .A(n10558), .B(n9637), .Y(n5305) );
  AOI22X1TS U11263 ( .A0(n11543), .A1(n11040), .B0(n12309), .B1(n12651), .Y(
        n2133) );
  AOI22X1TS U11264 ( .A0(n3756), .A1(n11721), .B0(n10477), .B1(n12509), .Y(
        n4653) );
  INVX2TS U11265 ( .A(n5593), .Y(n11716) );
  INVX2TS U11266 ( .A(n12330), .Y(n10014) );
  CLKBUFX2TS U11267 ( .A(n10398), .Y(n3724) );
  INVX1TS U11268 ( .A(n4480), .Y(n10803) );
  INVX1TS U11269 ( .A(n7130), .Y(n12090) );
  CLKINVX2TS U11270 ( .A(n10688), .Y(n9818) );
  INVX1TS U11271 ( .A(n5550), .Y(n12273) );
  INVX1TS U11272 ( .A(n3558), .Y(n12437) );
  CLKINVX2TS U11273 ( .A(n11370), .Y(n9916) );
  CLKINVX2TS U11274 ( .A(n7182), .Y(n11844) );
  INVX2TS U11275 ( .A(n3567), .Y(n10901) );
  INVX2TS U11276 ( .A(n7396), .Y(n10294) );
  CLKINVX2TS U11277 ( .A(n12059), .Y(n10481) );
  AOI22X1TS U11278 ( .A0(n11797), .A1(n12378), .B0(n10379), .B1(n11272), .Y(
        n4278) );
  CLKINVX2TS U11279 ( .A(n7169), .Y(n11469) );
  INVX1TS U11280 ( .A(n5550), .Y(n12271) );
  CLKINVX2TS U11281 ( .A(n10733), .Y(n12321) );
  INVX2TS U11282 ( .A(n5593), .Y(n11718) );
  INVX2TS U11283 ( .A(n2380), .Y(n11483) );
  INVX2TS U11284 ( .A(n4075), .Y(n9138) );
  CLKINVX2TS U11285 ( .A(n2687), .Y(n11435) );
  CLKINVX2TS U11286 ( .A(n12365), .Y(n9979) );
  AOI22X1TS U11287 ( .A0(n10586), .A1(n11712), .B0(n10441), .B1(n12521), .Y(
        n6453) );
  CLKINVX2TS U11288 ( .A(n2247), .Y(n10219) );
  INVX2TS U11289 ( .A(n3528), .Y(n10915) );
  INVX2TS U11290 ( .A(n2687), .Y(n11434) );
  CLKINVX2TS U11291 ( .A(n2559), .Y(n10176) );
  INVX2TS U11292 ( .A(n1819), .Y(n12360) );
  CLKINVX2TS U11293 ( .A(n3757), .Y(n10822) );
  INVX1TS U11294 ( .A(n3597), .Y(n12421) );
  CLKINVX2TS U11295 ( .A(n5512), .Y(n10919) );
  INVX2TS U11296 ( .A(n5908), .Y(n11012) );
  CLKINVX2TS U11297 ( .A(n11634), .Y(n10594) );
  CLKINVX2TS U11298 ( .A(n12652), .Y(n11859) );
  CLKINVX2TS U11299 ( .A(n12059), .Y(n10480) );
  INVX2TS U11300 ( .A(n1713), .Y(n11619) );
  CLKINVX2TS U11301 ( .A(n11635), .Y(n10595) );
  INVX2TS U11302 ( .A(n10782), .Y(n10147) );
  CLKINVX2TS U11303 ( .A(n11228), .Y(n10500) );
  INVX1TS U11304 ( .A(n5365), .Y(n10869) );
  CLKINVX2TS U11305 ( .A(n10840), .Y(n10989) );
  INVX1TS U11306 ( .A(n4108), .Y(n10779) );
  INVX2TS U11307 ( .A(n3895), .Y(n9655) );
  INVX1TS U11308 ( .A(n3528), .Y(n10917) );
  INVX2TS U11309 ( .A(n7076), .Y(n12456) );
  CLKINVX2TS U11310 ( .A(n2720), .Y(n11429) );
  INVX1TS U11311 ( .A(n4052), .Y(n10768) );
  INVX2TS U11312 ( .A(n3795), .Y(n12214) );
  INVX2TS U11313 ( .A(n5317), .Y(n9637) );
  INVX2TS U11314 ( .A(n12454), .Y(n9692) );
  INVX2TS U11315 ( .A(n1846), .Y(n10279) );
  CLKINVX2TS U11316 ( .A(n11463), .Y(n10038) );
  CLKINVX1TS U11317 ( .A(n2380), .Y(n11484) );
  INVX2TS U11318 ( .A(n5582), .Y(n10479) );
  INVX2TS U11319 ( .A(n7068), .Y(n11771) );
  CLKINVX2TS U11320 ( .A(n7163), .Y(n11818) );
  CLKBUFX2TS U11321 ( .A(n11311), .Y(n5527) );
  INVX1TS U11322 ( .A(n4108), .Y(n10780) );
  INVX2TS U11323 ( .A(n11368), .Y(n9915) );
  INVX1TS U11324 ( .A(n10626), .Y(n11010) );
  CLKINVX2TS U11325 ( .A(n7169), .Y(n11468) );
  INVX2TS U11326 ( .A(n12318), .Y(n9688) );
  INVX2TS U11327 ( .A(n3729), .Y(n12222) );
  INVX1TS U11328 ( .A(n6006), .Y(n11395) );
  CLKBUFX2TS U11329 ( .A(n11794), .Y(n7167) );
  INVX1TS U11330 ( .A(n5908), .Y(n11013) );
  INVX2TS U11331 ( .A(n3544), .Y(n12445) );
  INVX2TS U11332 ( .A(n2308), .Y(n10981) );
  INVX2TS U11333 ( .A(n5700), .Y(n9715) );
  CLKINVX2TS U11334 ( .A(n1844), .Y(n9992) );
  INVX2TS U11335 ( .A(n12643), .Y(n10357) );
  INVX2TS U11336 ( .A(n11654), .Y(n9822) );
  CLKINVX1TS U11337 ( .A(n2039), .Y(n11046) );
  INVX2TS U11338 ( .A(n11113), .Y(n11444) );
  INVX2TS U11339 ( .A(n2022), .Y(n10611) );
  CLKINVX2TS U11340 ( .A(n7122), .Y(n12464) );
  INVX2TS U11341 ( .A(n5725), .Y(n9719) );
  CLKINVX2TS U11342 ( .A(n2066), .Y(n10596) );
  INVX1TS U11343 ( .A(n5908), .Y(n11014) );
  INVX2TS U11344 ( .A(n12650), .Y(n11857) );
  INVX1TS U11345 ( .A(n5365), .Y(n10870) );
  CLKINVX2TS U11346 ( .A(n7241), .Y(n11487) );
  INVX2TS U11347 ( .A(n10624), .Y(n11009) );
  CLKINVX2TS U11348 ( .A(n2039), .Y(n11047) );
  INVX2TS U11349 ( .A(n7607), .Y(n11908) );
  INVX2TS U11350 ( .A(n11654), .Y(n9821) );
  CLKINVX2TS U11351 ( .A(n5512), .Y(n10918) );
  INVX2TS U11352 ( .A(n7975), .Y(n12597) );
  INVX2TS U11353 ( .A(n7591), .Y(n12178) );
  CLKINVX2TS U11354 ( .A(n10986), .Y(n11882) );
  INVX1TS U11355 ( .A(n2483), .Y(n10519) );
  CLKBUFX2TS U11356 ( .A(n10021), .Y(n7893) );
  CLKINVX2TS U11357 ( .A(n10735), .Y(n12319) );
  CLKBUFX2TS U11358 ( .A(n11198), .Y(n7629) );
  INVX2TS U11359 ( .A(n5326), .Y(n10853) );
  INVX2TS U11360 ( .A(n7607), .Y(n11909) );
  CLKINVX1TS U11361 ( .A(n12570), .Y(n9641) );
  CLKINVX2TS U11362 ( .A(n8193), .Y(n11188) );
  CLKINVX2TS U11363 ( .A(n12324), .Y(n10694) );
  CLKINVX2TS U11364 ( .A(n1693), .Y(n11636) );
  INVX2TS U11365 ( .A(n7975), .Y(n12596) );
  INVX1TS U11366 ( .A(n11114), .Y(n11445) );
  INVX2TS U11367 ( .A(n3870), .Y(n9659) );
  INVX1TS U11368 ( .A(n2032), .Y(n12092) );
  INVX2TS U11369 ( .A(n1989), .Y(n10619) );
  CLKINVX2TS U11370 ( .A(n8193), .Y(n11187) );
  INVX2TS U11371 ( .A(n12193), .Y(n10287) );
  INVX1TS U11372 ( .A(n11021), .Y(n11023) );
  INVX2TS U11373 ( .A(n7105), .Y(n10253) );
  CLKINVX2TS U11374 ( .A(n1803), .Y(n12161) );
  INVX2TS U11375 ( .A(n11021), .Y(n11022) );
  INVX1TS U11376 ( .A(n2069), .Y(n11041) );
  CLKBUFX2TS U11377 ( .A(n10053), .Y(n7231) );
  INVX2TS U11378 ( .A(n2032), .Y(n12091) );
  INVX2TS U11379 ( .A(n12622), .Y(n10187) );
  CLKBUFX2TS U11380 ( .A(n11290), .Y(n3772) );
  CLKINVX2TS U11381 ( .A(n11130), .Y(n11120) );
  INVX2TS U11382 ( .A(n11459), .Y(n9956) );
  INVX2TS U11383 ( .A(n2559), .Y(n10175) );
  INVX2TS U11384 ( .A(n2168), .Y(n10587) );
  INVX2TS U11385 ( .A(n11440), .Y(n10191) );
  CLKINVX2TS U11386 ( .A(n5388), .Y(n10452) );
  INVX2TS U11387 ( .A(n11089), .Y(n10252) );
  INVX1TS U11388 ( .A(n3795), .Y(n12216) );
  INVX2TS U11389 ( .A(n12653), .Y(n11858) );
  INVX1TS U11390 ( .A(n11021), .Y(n11024) );
  INVX1TS U11391 ( .A(n2168), .Y(n10588) );
  INVX2TS U11392 ( .A(n2720), .Y(n11428) );
  INVX2TS U11393 ( .A(n10965), .Y(n10966) );
  INVX2TS U11394 ( .A(n2247), .Y(n10220) );
  INVX2TS U11395 ( .A(n5381), .Y(n12399) );
  CLKINVX2TS U11396 ( .A(n2066), .Y(n10598) );
  CLKINVX2TS U11397 ( .A(n11442), .Y(n10192) );
  INVX2TS U11398 ( .A(n2650), .Y(n9923) );
  INVX2TS U11399 ( .A(n7607), .Y(n11910) );
  CLKINVX2TS U11400 ( .A(n1989), .Y(n10620) );
  CLKBUFX2TS U11401 ( .A(n11170), .Y(n7276) );
  INVX2TS U11402 ( .A(n2039), .Y(n11045) );
  CLKINVX2TS U11403 ( .A(n11283), .Y(n9950) );
  INVX2TS U11404 ( .A(n1960), .Y(n12110) );
  INVX2TS U11405 ( .A(n7285), .Y(n11091) );
  INVX1TS U11406 ( .A(n5550), .Y(n12274) );
  INVX2TS U11407 ( .A(n11281), .Y(n9949) );
  INVX2TS U11408 ( .A(n11520), .Y(n10304) );
  INVX1TS U11409 ( .A(n2168), .Y(n10589) );
  INVX1TS U11410 ( .A(n7591), .Y(n12179) );
  INVX2TS U11411 ( .A(n1909), .Y(n10255) );
  CLKINVX2TS U11412 ( .A(n1693), .Y(n11638) );
  CLKINVX2TS U11413 ( .A(n12058), .Y(n10482) );
  CLKINVX1TS U11414 ( .A(n5342), .Y(n12384) );
  CLKINVX2TS U11415 ( .A(n10799), .Y(n10943) );
  INVX1TS U11416 ( .A(n3729), .Y(n12221) );
  CLKINVX2TS U11417 ( .A(n11105), .Y(n10276) );
  INVX2TS U11418 ( .A(n10988), .Y(n11883) );
  CLKINVX2TS U11419 ( .A(n11154), .Y(n11142) );
  INVX1TS U11420 ( .A(n4052), .Y(n10767) );
  INVX2TS U11421 ( .A(n7259), .Y(n9471) );
  INVX2TS U11422 ( .A(n10882), .Y(n10787) );
  CLKINVX2TS U11423 ( .A(n12326), .Y(n10693) );
  CLKINVX2TS U11424 ( .A(n7539), .Y(n10678) );
  CLKINVX2TS U11425 ( .A(n2590), .Y(n10956) );
  CLKINVX2TS U11426 ( .A(n3757), .Y(n10823) );
  INVX2TS U11427 ( .A(n11506), .Y(n10292) );
  CLKINVX2TS U11428 ( .A(n5388), .Y(n10453) );
  INVX2TS U11429 ( .A(n4108), .Y(n10778) );
  INVX2TS U11430 ( .A(n12367), .Y(n9980) );
  INVX1TS U11431 ( .A(n5395), .Y(n12409) );
  INVX2TS U11432 ( .A(n4052), .Y(n10766) );
  CLKINVX2TS U11433 ( .A(n3691), .Y(n10849) );
  CLKINVX2TS U11434 ( .A(n1803), .Y(n12159) );
  CLKINVX2TS U11435 ( .A(n2424), .Y(n11470) );
  INVX2TS U11436 ( .A(n2590), .Y(n10954) );
  INVX1TS U11437 ( .A(n4239), .Y(n11218) );
  CLKINVX2TS U11438 ( .A(n10637), .Y(n10998) );
  INVX1TS U11439 ( .A(n3528), .Y(n10916) );
  INVX2TS U11440 ( .A(n11106), .Y(n10275) );
  INVX2TS U11441 ( .A(n5365), .Y(n10868) );
  CLKINVX2TS U11442 ( .A(n1713), .Y(n11618) );
  CLKBUFX2TS U11443 ( .A(n11338), .Y(n3706) );
  INVX1TS U11444 ( .A(n1713), .Y(n11620) );
  CLKINVX2TS U11445 ( .A(n3757), .Y(n10821) );
  INVX2TS U11446 ( .A(n7241), .Y(n11485) );
  AOI22X1TS U11447 ( .A0(n5445), .A1(n11694), .B0(n10423), .B1(n12505), .Y(
        n6381) );
  INVX2TS U11448 ( .A(n3519), .Y(n9634) );
  INVX2TS U11449 ( .A(n1803), .Y(n12160) );
  INVX2TS U11450 ( .A(n11112), .Y(n11443) );
  CLKBUFX2TS U11451 ( .A(n11953), .Y(n2041) );
  INVX2TS U11452 ( .A(n5931), .Y(n9349) );
  AOI22X1TS U11453 ( .A0(n3690), .A1(n11739), .B0(n10495), .B1(n12525), .Y(
        n4581) );
  INVX2TS U11454 ( .A(n10972), .Y(n11907) );
  INVX1TS U11455 ( .A(n1960), .Y(n12112) );
  INVX2TS U11456 ( .A(n11152), .Y(n11141) );
  INVX2TS U11457 ( .A(n5381), .Y(n12401) );
  CLKINVX2TS U11458 ( .A(n7539), .Y(n10677) );
  CLKBUFX2TS U11459 ( .A(n11642), .Y(n1691) );
  CLKINVX2TS U11460 ( .A(n7122), .Y(n12465) );
  INVX2TS U11461 ( .A(n12193), .Y(n10288) );
  CLKINVX2TS U11462 ( .A(n1675), .Y(n12562) );
  CLKINVX2TS U11463 ( .A(n5512), .Y(n10920) );
  AOI22X1TS U11464 ( .A0(n12278), .A1(n12537), .B0(n11740), .B1(n5962), .Y(
        n6342) );
  INVX1TS U11465 ( .A(n5381), .Y(n12400) );
  INVX2TS U11466 ( .A(n1675), .Y(n12565) );
  INVX1TS U11467 ( .A(n7130), .Y(n12089) );
  INVX2TS U11468 ( .A(n5550), .Y(n12272) );
  INVX2TS U11469 ( .A(n7550), .Y(n10328) );
  INVX2TS U11470 ( .A(n2069), .Y(n11040) );
  CLKINVX1TS U11471 ( .A(n1989), .Y(n10621) );
  CLKINVX2TS U11472 ( .A(n12624), .Y(n10188) );
  INVX1TS U11473 ( .A(n3567), .Y(n10900) );
  INVX2TS U11474 ( .A(n2066), .Y(n10597) );
  CLKINVX2TS U11475 ( .A(n2590), .Y(n10955) );
  CLKINVX2TS U11476 ( .A(n11132), .Y(n11121) );
  INVX1TS U11477 ( .A(n10965), .Y(n10967) );
  INVX2TS U11478 ( .A(n7285), .Y(n11093) );
  CLKINVX1TS U11479 ( .A(n2424), .Y(n11472) );
  INVX1TS U11480 ( .A(n2032), .Y(n12093) );
  CLKINVX2TS U11481 ( .A(n10635), .Y(n10997) );
  INVX2TS U11482 ( .A(n12451), .Y(n9693) );
  INVX2TS U11483 ( .A(n11460), .Y(n9955) );
  INVX2TS U11484 ( .A(n12315), .Y(n9689) );
  INVX2TS U11485 ( .A(n12046), .Y(n9908) );
  INVX2TS U11486 ( .A(n1693), .Y(n11637) );
  CLKINVX2TS U11487 ( .A(n11629), .Y(n10608) );
  INVX1TS U11488 ( .A(n1960), .Y(n12111) );
  CLKINVX2TS U11489 ( .A(n11089), .Y(n10251) );
  INVX2TS U11490 ( .A(n1751), .Y(n11601) );
  CLKINVX2TS U11491 ( .A(n2308), .Y(n10982) );
  INVX1TS U11492 ( .A(n9766), .Y(n11981) );
  INVX2TS U11493 ( .A(n10397), .Y(n9901) );
  INVX2TS U11494 ( .A(n7739), .Y(n11926) );
  CLKINVX2TS U11495 ( .A(n10927), .Y(n10755) );
  CLKBUFX2TS U11496 ( .A(n10073), .Y(n7827) );
  INVX1TS U11497 ( .A(n7322), .Y(n12142) );
  CLKINVX2TS U11498 ( .A(n5299), .Y(n12204) );
  CLKINVX2TS U11499 ( .A(n11376), .Y(n10407) );
  INVX1TS U11500 ( .A(n5579), .Y(n11330) );
  CLKINVX2TS U11501 ( .A(n10798), .Y(n9922) );
  CLKINVX2TS U11502 ( .A(n6015), .Y(n11402) );
  INVX2TS U11503 ( .A(n5484), .Y(n12264) );
  INVX2TS U11504 ( .A(n6006), .Y(n11396) );
  INVX2TS U11505 ( .A(n7846), .Y(n11615) );
  INVX2TS U11506 ( .A(n5579), .Y(n11331) );
  INVX1TS U11507 ( .A(n7322), .Y(n12143) );
  CLKINVX2TS U11508 ( .A(n10786), .Y(n11708) );
  CLKINVX2TS U11509 ( .A(n5342), .Y(n12385) );
  CLKINVX2TS U11510 ( .A(n3501), .Y(n12283) );
  INVX2TS U11511 ( .A(n3795), .Y(n12213) );
  CLKINVX2TS U11512 ( .A(n11343), .Y(n9966) );
  CLKINVX2TS U11513 ( .A(n10841), .Y(n10990) );
  CLKINVX2TS U11514 ( .A(n3516), .Y(n10498) );
  INVX2TS U11515 ( .A(n5875), .Y(n9334) );
  INVX2TS U11516 ( .A(n5326), .Y(n10851) );
  INVX2TS U11517 ( .A(n7495), .Y(n11558) );
  CLKINVX2TS U11518 ( .A(n5293), .Y(n10825) );
  INVX2TS U11519 ( .A(n7105), .Y(n10254) );
  CLKINVX2TS U11520 ( .A(n3996), .Y(n10402) );
  INVX2TS U11521 ( .A(n10951), .Y(n10819) );
  INVX2TS U11522 ( .A(n10801), .Y(n10944) );
  CLKBUFX2TS U11523 ( .A(n10525), .Y(n5479) );
  INVX2TS U11524 ( .A(n7739), .Y(n11927) );
  INVX1TS U11525 ( .A(n6296), .Y(n12299) );
  INVX1TS U11526 ( .A(n3795), .Y(n12215) );
  CLKINVX1TS U11527 ( .A(n10953), .Y(n10820) );
  CLKINVX2TS U11528 ( .A(n3583), .Y(n12430) );
  INVX2TS U11529 ( .A(n4239), .Y(n11220) );
  INVX2TS U11530 ( .A(n5593), .Y(n11717) );
  CLKINVX2TS U11531 ( .A(n12017), .Y(n9675) );
  CLKINVX2TS U11532 ( .A(n5349), .Y(n10436) );
  INVX2TS U11533 ( .A(n5428), .Y(n11976) );
  INVX2TS U11534 ( .A(n5578), .Y(n10177) );
  INVX2TS U11535 ( .A(n7259), .Y(n9472) );
  INVX1TS U11536 ( .A(n5356), .Y(n12393) );
  AOI22X1TS U11537 ( .A0(n10584), .A1(n11453), .B0(n10231), .B1(n1820), .Y(
        n3097) );
  INVX2TS U11538 ( .A(n4259), .Y(n10125) );
  AOI22X1TS U11539 ( .A0(n11797), .A1(n12594), .B0(n10380), .B1(n3992), .Y(
        n4352) );
  CLKINVX2TS U11540 ( .A(n4350), .Y(n9661) );
  INVX2TS U11541 ( .A(n7130), .Y(n12088) );
  CLKINVX2TS U11542 ( .A(n11322), .Y(n9912) );
  INVX1TS U11543 ( .A(n5972), .Y(n12294) );
  INVX1TS U11544 ( .A(n5484), .Y(n12263) );
  INVX1TS U11545 ( .A(n7076), .Y(n12455) );
  INVX2TS U11546 ( .A(n4351), .Y(n9665) );
  INVX1TS U11547 ( .A(n5852), .Y(n11001) );
  CLKINVX2TS U11548 ( .A(n12621), .Y(n10144) );
  INVX2TS U11549 ( .A(n6296), .Y(n12298) );
  CLKINVX2TS U11550 ( .A(n12043), .Y(n9907) );
  CLKBUFX2TS U11551 ( .A(n11597), .Y(n7651) );
  CLKINVX2TS U11552 ( .A(n3648), .Y(n10872) );
  CLKINVX2TS U11553 ( .A(n7495), .Y(n11557) );
  CLKINVX1TS U11554 ( .A(n10800), .Y(n10945) );
  CLKINVX2TS U11555 ( .A(n10971), .Y(n11905) );
  CLKINVX1TS U11556 ( .A(n2650), .Y(n9924) );
  INVX2TS U11557 ( .A(n10771), .Y(n10391) );
  INVX2TS U11558 ( .A(n6026), .Y(n10242) );
  INVX2TS U11559 ( .A(n11439), .Y(n10590) );
  INVX2TS U11560 ( .A(n7739), .Y(n11928) );
  INVX1TS U11561 ( .A(n5484), .Y(n12266) );
  CLKINVX2TS U11562 ( .A(n9998), .Y(n10413) );
  INVX2TS U11563 ( .A(n11233), .Y(n9945) );
  CLKINVX2TS U11564 ( .A(n10842), .Y(n10991) );
  CLKINVX2TS U11565 ( .A(n11235), .Y(n9946) );
  INVX2TS U11566 ( .A(n6153), .Y(n9758) );
  INVX2TS U11567 ( .A(n6010), .Y(n9989) );
  INVX2TS U11568 ( .A(n12620), .Y(n10143) );
  INVX2TS U11569 ( .A(n6287), .Y(n10249) );
  INVX1TS U11570 ( .A(n6010), .Y(n9990) );
  INVX2TS U11571 ( .A(n5972), .Y(n12292) );
  INVX1TS U11572 ( .A(n5299), .Y(n12205) );
  INVX2TS U11573 ( .A(n6015), .Y(n11401) );
  INVX2TS U11574 ( .A(n10655), .Y(n10315) );
  INVX2TS U11575 ( .A(n10796), .Y(n9921) );
  INVX2TS U11576 ( .A(n11342), .Y(n9965) );
  CLKINVX2TS U11577 ( .A(n10952), .Y(n10818) );
  INVX2TS U11578 ( .A(n5299), .Y(n12203) );
  CLKINVX1TS U11579 ( .A(n3590), .Y(n10463) );
  INVX2TS U11580 ( .A(n4131), .Y(n9150) );
  CLKINVX2TS U11581 ( .A(n5349), .Y(n10435) );
  INVX1TS U11582 ( .A(n5972), .Y(n12293) );
  INVX1TS U11583 ( .A(n10769), .Y(n10390) );
  CLKBUFX2TS U11584 ( .A(n10562), .Y(n5316) );
  INVX1TS U11585 ( .A(n7076), .Y(n12457) );
  CLKINVX1TS U11586 ( .A(n7495), .Y(n11559) );
  CLKINVX2TS U11587 ( .A(n11153), .Y(n11143) );
  CLKINVX2TS U11588 ( .A(n11376), .Y(n10406) );
  INVX2TS U11589 ( .A(n6154), .Y(n9763) );
  CLKINVX2TS U11590 ( .A(n3583), .Y(n12427) );
  INVX2TS U11591 ( .A(n3954), .Y(n10148) );
  CLKINVX2TS U11592 ( .A(n6154), .Y(n9762) );
  INVX2TS U11593 ( .A(n6287), .Y(n10250) );
  INVX2TS U11594 ( .A(n5800), .Y(n10522) );
  CLKINVX2TS U11595 ( .A(n6153), .Y(n9759) );
  INVX2TS U11596 ( .A(n6026), .Y(n10241) );
  INVX2TS U11597 ( .A(n3567), .Y(n10899) );
  CLKINVX2TS U11598 ( .A(n5428), .Y(n11977) );
  INVX2TS U11599 ( .A(n10655), .Y(n10316) );
  CLKBUFX2TS U11600 ( .A(n10554), .Y(n5298) );
  INVX2TS U11601 ( .A(n9766), .Y(n11979) );
  INVX2TS U11602 ( .A(n12570), .Y(n9640) );
  INVX2TS U11603 ( .A(n6006), .Y(n11397) );
  INVX1TS U11604 ( .A(n4492), .Y(n9190) );
  INVX1TS U11605 ( .A(n7655), .Y(n12184) );
  CLKINVX2TS U11606 ( .A(n12071), .Y(n10502) );
  CLKBUFX2TS U11607 ( .A(n11741), .Y(n5600) );
  CLKINVX2TS U11608 ( .A(n5800), .Y(n10521) );
  CLKINVX2TS U11609 ( .A(n10882), .Y(n10789) );
  INVX1TS U11610 ( .A(n2483), .Y(n10520) );
  CLKINVX2TS U11611 ( .A(n1720), .Y(n10667) );
  CLKINVX2TS U11612 ( .A(n3516), .Y(n10499) );
  INVX1TS U11613 ( .A(n6296), .Y(n12300) );
  INVX2TS U11614 ( .A(n11320), .Y(n9911) );
  INVX1TS U11615 ( .A(n9767), .Y(n11980) );
  INVX1TS U11616 ( .A(n5852), .Y(n11002) );
  NOR2X1TS U11617 ( .A(n11957), .B(n11145), .Y(n7659) );
  AOI22X1TS U11618 ( .A0(n11683), .A1(n12576), .B0(n10563), .B1(n5785), .Y(
        n6155) );
  CLKINVX2TS U11619 ( .A(n5314), .Y(n10416) );
  INVX2TS U11620 ( .A(n5415), .Y(n10154) );
  INVX1TS U11621 ( .A(n3501), .Y(n12284) );
  INVX2TS U11622 ( .A(n5582), .Y(n10478) );
  INVX1TS U11623 ( .A(n5326), .Y(n10852) );
  CLKINVX2TS U11624 ( .A(n1751), .Y(n11602) );
  INVX2TS U11625 ( .A(n12328), .Y(n10013) );
  CLKINVX2TS U11626 ( .A(n3648), .Y(n10871) );
  INVX2TS U11627 ( .A(n4480), .Y(n10802) );
  INVX2TS U11628 ( .A(n5579), .Y(n11329) );
  INVX2TS U11629 ( .A(n4239), .Y(n11219) );
  INVX2TS U11630 ( .A(n2424), .Y(n11471) );
  INVX1TS U11631 ( .A(n7322), .Y(n12141) );
  INVX2TS U11632 ( .A(n10785), .Y(n11707) );
  INVX2TS U11633 ( .A(n11268), .Y(n9913) );
  INVX2TS U11634 ( .A(n11437), .Y(n10591) );
  INVX1TS U11635 ( .A(n2022), .Y(n10610) );
  INVX1TS U11636 ( .A(n4243), .Y(n9934) );
  INVX1TS U11637 ( .A(n10883), .Y(n10788) );
  CLKINVX2TS U11638 ( .A(n7122), .Y(n12463) );
  INVX2TS U11639 ( .A(n5578), .Y(n10178) );
  CLKBUFX2TS U11640 ( .A(n11860), .Y(n7734) );
  CLKBUFX2TS U11641 ( .A(n10379), .Y(n3518) );
  INVX2TS U11642 ( .A(n7068), .Y(n11770) );
  INVX2TS U11643 ( .A(n7655), .Y(n12185) );
  CLKBUFX2TS U11644 ( .A(n12486), .Y(n7314) );
  INVX2TS U11645 ( .A(n7682), .Y(n10066) );
  CLKINVX2TS U11646 ( .A(n10973), .Y(n11906) );
  CLKINVX2TS U11647 ( .A(n7682), .Y(n10065) );
  CLKINVX2TS U11648 ( .A(n10733), .Y(n12320) );
  CLKINVX2TS U11649 ( .A(n12599), .Y(n10211) );
  CLKINVX2TS U11650 ( .A(n10928), .Y(n10756) );
  INVX2TS U11651 ( .A(n9632), .Y(n10212) );
  CLKINVX2TS U11652 ( .A(n10987), .Y(n11881) );
  INVX2TS U11653 ( .A(n4492), .Y(n9189) );
  INVX2TS U11654 ( .A(n5852), .Y(n11000) );
  CLKINVX2TS U11655 ( .A(n7182), .Y(n11843) );
  INVX1TS U11656 ( .A(n5875), .Y(n9335) );
  INVX1TS U11657 ( .A(n7655), .Y(n12183) );
  INVX2TS U11658 ( .A(n4259), .Y(n10126) );
  CLKINVX2TS U11659 ( .A(n7068), .Y(n11772) );
  CLKINVX2TS U11660 ( .A(n10397), .Y(n9902) );
  INVX2TS U11661 ( .A(n1844), .Y(n9991) );
  INVX2TS U11662 ( .A(n4243), .Y(n9933) );
  CLKINVX2TS U11663 ( .A(n3590), .Y(n10464) );
  INVX2TS U11664 ( .A(n7846), .Y(n11616) );
  INVX2TS U11665 ( .A(n11461), .Y(n10037) );
  INVX2TS U11666 ( .A(n4350), .Y(n9660) );
  CLKBUFX2TS U11667 ( .A(n10369), .Y(n3500) );
  CLKINVX2TS U11668 ( .A(n5446), .Y(n10891) );
  INVX2TS U11669 ( .A(n7550), .Y(n10329) );
  CLKINVX2TS U11670 ( .A(n1758), .Y(n10653) );
  CLKINVX2TS U11671 ( .A(n7241), .Y(n11486) );
  INVX2TS U11672 ( .A(n7846), .Y(n11617) );
  CLKINVX2TS U11673 ( .A(n10784), .Y(n11709) );
  CLKINVX2TS U11674 ( .A(n11267), .Y(n9914) );
  CLKINVX2TS U11675 ( .A(n4351), .Y(n9664) );
  CLKBUFX2TS U11676 ( .A(n11263), .Y(n5461) );
  CLKBUFX2TS U11677 ( .A(n10429), .Y(n3991) );
  CLKBUFX2TS U11678 ( .A(n10337), .Y(n7815) );
  OR2X2TS U11679 ( .A(n9873), .B(n7489), .Y(n7666) );
  INVX2TS U11680 ( .A(n1692), .Y(n11642) );
  INVX2TS U11681 ( .A(n7715), .Y(n9861) );
  INVX2TS U11682 ( .A(n7716), .Y(n10073) );
  INVX2TS U11683 ( .A(n3692), .Y(n12404) );
  INVX1TS U11684 ( .A(n3738), .Y(n12514) );
  INVX2TS U11685 ( .A(n2256), .Y(n9947) );
  INVX2TS U11686 ( .A(n9626), .Y(n9627) );
  CLKBUFX2TS U11687 ( .A(n10235), .Y(n2145) );
  INVX2TS U11688 ( .A(n10376), .Y(n10136) );
  CLKINVX2TS U11689 ( .A(n5544), .Y(n11312) );
  INVX2TS U11690 ( .A(n7512), .Y(n11563) );
  CLKINVX1TS U11691 ( .A(n5445), .Y(n10461) );
  CLKBUFX2TS U11692 ( .A(n9729), .Y(n1714) );
  INVX2TS U11693 ( .A(n5328), .Y(n10421) );
  INVX1TS U11694 ( .A(n7141), .Y(n11457) );
  CLKINVX2TS U11695 ( .A(n3956), .Y(n11715) );
  INVX1TS U11696 ( .A(n7253), .Y(n10022) );
  CLKINVX2TS U11697 ( .A(n7668), .Y(n11598) );
  INVX1TS U11698 ( .A(n5559), .Y(n12526) );
  INVX1TS U11699 ( .A(n7695), .Y(n11145) );
  INVX2TS U11700 ( .A(n5493), .Y(n12511) );
  INVX2TS U11701 ( .A(n12082), .Y(n10025) );
  INVX2TS U11702 ( .A(n3738), .Y(n12517) );
  INVX2TS U11703 ( .A(n7526), .Y(n10053) );
  INVX2TS U11704 ( .A(n4501), .Y(n10813) );
  CLKINVX2TS U11705 ( .A(n3690), .Y(n10446) );
  INVX2TS U11706 ( .A(n5513), .Y(n12424) );
  INVX1TS U11707 ( .A(n10681), .Y(n11078) );
  INVX2TS U11708 ( .A(n6039), .Y(n10562) );
  INVX2TS U11709 ( .A(n3569), .Y(n10475) );
  INVX2TS U11710 ( .A(n1822), .Y(n11912) );
  CLKINVX2TS U11711 ( .A(n1676), .Y(n9765) );
  INVX2TS U11712 ( .A(n3643), .Y(n12030) );
  INVX2TS U11713 ( .A(n1810), .Y(n11588) );
  CLKBUFX2TS U11714 ( .A(n11815), .Y(n2466) );
  INVX2TS U11715 ( .A(n6012), .Y(n10554) );
  CLKBUFX2TS U11716 ( .A(n10565), .Y(n1740) );
  INVX1TS U11717 ( .A(n11026), .Y(n11605) );
  INVX2TS U11718 ( .A(n7131), .Y(n12094) );
  CLKBUFX2TS U11719 ( .A(n12575), .Y(n5296) );
  INVX2TS U11720 ( .A(n4245), .Y(n10369) );
  INVX2TS U11721 ( .A(n5743), .Y(n11740) );
  OR2X2TS U11722 ( .A(n9951), .B(n2508), .Y(n2629) );
  INVX1TS U11723 ( .A(n10719), .Y(n11124) );
  CLKBUFX2TS U11724 ( .A(n12593), .Y(n3498) );
  INVX1TS U11725 ( .A(n3738), .Y(n12515) );
  CLKBUFX2TS U11726 ( .A(n10111), .Y(n3912) );
  INVX2TS U11727 ( .A(n4272), .Y(n10379) );
  INVX2TS U11728 ( .A(n10371), .Y(n10128) );
  INVX2TS U11729 ( .A(n7393), .Y(n11886) );
  INVX1TS U11730 ( .A(n3804), .Y(n12499) );
  CLKBUFX2TS U11731 ( .A(n9987), .Y(n1875) );
  CLKBUFX2TS U11732 ( .A(n10197), .Y(n5671) );
  CLKINVX1TS U11733 ( .A(n4113), .Y(n10389) );
  INVX2TS U11734 ( .A(n2020), .Y(n12333) );
  AND2X2TS U11735 ( .A(n4925), .B(n4903), .Y(n3827) );
  OR2X2TS U11736 ( .A(n8022), .B(n9873), .Y(n7476) );
  INVX2TS U11737 ( .A(n7393), .Y(n11884) );
  INVX2TS U11738 ( .A(n10717), .Y(n11123) );
  AND2X2TS U11739 ( .A(n4903), .B(n3830), .Y(n4013) );
  CLKINVX2TS U11740 ( .A(n3758), .Y(n12395) );
  CLKBUFX2TS U11741 ( .A(n10195), .Y(n2171) );
  INVX1TS U11742 ( .A(n4272), .Y(n10380) );
  INVX2TS U11743 ( .A(n10795), .Y(n10160) );
  CLKINVX2TS U11744 ( .A(n11798), .Y(n9169) );
  CLKBUFX2TS U11745 ( .A(n9740), .Y(n1749) );
  CLKBUFX2TS U11746 ( .A(n11920), .Y(n7310) );
  INVX2TS U11747 ( .A(n7662), .Y(n12488) );
  INVX2TS U11748 ( .A(n1676), .Y(n9764) );
  INVX2TS U11749 ( .A(n5511), .Y(n10470) );
  INVX1TS U11750 ( .A(n7662), .Y(n12489) );
  INVX2TS U11751 ( .A(n7331), .Y(n11860) );
  INVX2TS U11752 ( .A(n10371), .Y(n10127) );
  INVX2TS U11753 ( .A(n3956), .Y(n11713) );
  INVX2TS U11754 ( .A(n7486), .Y(n12632) );
  INVX2TS U11755 ( .A(n4057), .Y(n10398) );
  CLKINVX1TS U11756 ( .A(n5913), .Y(n10536) );
  INVX2TS U11757 ( .A(n4113), .Y(n10387) );
  INVX1TS U11758 ( .A(n3643), .Y(n12032) );
  CLKBUFX2TS U11759 ( .A(n9930), .Y(n3490) );
  CLKINVX1TS U11760 ( .A(n7716), .Y(n10074) );
  CLKBUFX2TS U11761 ( .A(n10239), .Y(n2245) );
  CLKBUFX2TS U11762 ( .A(n12040), .Y(n5514) );
  INVX2TS U11763 ( .A(n7668), .Y(n11597) );
  INVX2TS U11764 ( .A(n5559), .Y(n12529) );
  INVX2TS U11765 ( .A(n7649), .Y(n12355) );
  INVX1TS U11766 ( .A(n4245), .Y(n10370) );
  INVX2TS U11767 ( .A(n5559), .Y(n12527) );
  INVX2TS U11768 ( .A(n3804), .Y(n12498) );
  INVX2TS U11769 ( .A(n7512), .Y(n11564) );
  INVX2TS U11770 ( .A(n7486), .Y(n12633) );
  INVX1TS U11771 ( .A(n1669), .Y(n11955) );
  INVX2TS U11772 ( .A(n10376), .Y(n10135) );
  INVX2TS U11773 ( .A(n11476), .Y(n9983) );
  INVX2TS U11774 ( .A(n2256), .Y(n9948) );
  INVX2TS U11775 ( .A(n7662), .Y(n12486) );
  INVX2TS U11776 ( .A(n3738), .Y(n12516) );
  CLKINVX1TS U11777 ( .A(n7438), .Y(n9501) );
  CLKBUFX2TS U11778 ( .A(n11509), .Y(n7693) );
  CLKBUFX2TS U11779 ( .A(n10539), .Y(n1702) );
  INVX2TS U11780 ( .A(n10793), .Y(n10159) );
  CLKBUFX2TS U11781 ( .A(n11536), .Y(n1974) );
  INVX2TS U11782 ( .A(n11855), .Y(n9520) );
  INVX2TS U11783 ( .A(n7073), .Y(n11432) );
  CLKBUFX2TS U11784 ( .A(n10285), .Y(n7737) );
  CLKINVX2TS U11785 ( .A(n1692), .Y(n11643) );
  INVX2TS U11786 ( .A(n7695), .Y(n11144) );
  CLKBUFX2TS U11787 ( .A(n9725), .Y(n1752) );
  INVX1TS U11788 ( .A(n3643), .Y(n12029) );
  INVX2TS U11789 ( .A(n3667), .Y(n12541) );
  INVX2TS U11790 ( .A(n11532), .Y(n10223) );
  INVX2TS U11791 ( .A(n7090), .Y(n11794) );
  INVX2TS U11792 ( .A(n3804), .Y(n12500) );
  INVX2TS U11793 ( .A(n5857), .Y(n10525) );
  CLKBUFX2TS U11794 ( .A(n10005), .Y(n7233) );
  CLKINVX2TS U11795 ( .A(n7649), .Y(n12357) );
  CLKINVX2TS U11796 ( .A(n11135), .Y(n11582) );
  INVX2TS U11797 ( .A(n5447), .Y(n12416) );
  INVX2TS U11798 ( .A(n3723), .Y(n11338) );
  INVX2TS U11799 ( .A(n7438), .Y(n9500) );
  INVX2TS U11800 ( .A(n7127), .Y(n11038) );
  INVX2TS U11801 ( .A(n11137), .Y(n11583) );
  CLKBUFX2TS U11802 ( .A(n10560), .Y(n1755) );
  CLKINVX2TS U11803 ( .A(n3667), .Y(n12539) );
  INVX2TS U11804 ( .A(n10599), .Y(n10289) );
  INVX2TS U11805 ( .A(n2323), .Y(n9944) );
  INVX2TS U11806 ( .A(n5493), .Y(n12513) );
  INVX2TS U11807 ( .A(n5367), .Y(n10439) );
  INVX1TS U11808 ( .A(n10962), .Y(n11544) );
  INVX2TS U11809 ( .A(n3690), .Y(n10447) );
  INVX2TS U11810 ( .A(n11466), .Y(n9971) );
  CLKBUFX2TS U11811 ( .A(n10459), .Y(n3671) );
  CLKBUFX2TS U11812 ( .A(n10874), .Y(n5506) );
  CLKINVX2TS U11813 ( .A(n3756), .Y(n10437) );
  CLKINVX2TS U11814 ( .A(n7077), .Y(n11778) );
  CLKBUFX2TS U11815 ( .A(n10015), .Y(n1811) );
  CLKINVX2TS U11816 ( .A(n5513), .Y(n12423) );
  INVX2TS U11817 ( .A(n1669), .Y(n11953) );
  INVX2TS U11818 ( .A(n3530), .Y(n10493) );
  CLKINVX2TS U11819 ( .A(n7090), .Y(n11796) );
  INVX2TS U11820 ( .A(n7141), .Y(n11455) );
  INVX2TS U11821 ( .A(n7127), .Y(n11037) );
  INVX1TS U11822 ( .A(n3804), .Y(n12501) );
  INVX2TS U11823 ( .A(n7238), .Y(n10622) );
  INVX2TS U11824 ( .A(n10599), .Y(n10290) );
  INVX2TS U11825 ( .A(n11466), .Y(n9972) );
  CLKBUFX2TS U11826 ( .A(n10263), .Y(n2312) );
  CLKBUFX2TS U11827 ( .A(n9975), .Y(n1938) );
  INVX2TS U11828 ( .A(n7077), .Y(n11776) );
  INVX2TS U11829 ( .A(n7393), .Y(n11885) );
  CLKBUFX2TS U11830 ( .A(n10911), .Y(n3685) );
  CLKBUFX2TS U11831 ( .A(n11209), .Y(n5844) );
  INVX2TS U11832 ( .A(n10961), .Y(n11543) );
  INVX1TS U11833 ( .A(n4113), .Y(n10388) );
  CLKBUFX2TS U11834 ( .A(n11392), .Y(n4100) );
  CLKINVX2TS U11835 ( .A(n11115), .Y(n11571) );
  CLKBUFX2TS U11836 ( .A(n10248), .Y(n2291) );
  INVX1TS U11837 ( .A(n7186), .Y(n11061) );
  CLKINVX2TS U11838 ( .A(n5447), .Y(n12415) );
  INVX2TS U11839 ( .A(n5345), .Y(n9635) );
  INVX1TS U11840 ( .A(n5559), .Y(n12528) );
  CLKBUFX2TS U11841 ( .A(n12149), .Y(n7185) );
  CLKINVX2TS U11842 ( .A(n4321), .Y(n12491) );
  CLKBUFX2TS U11843 ( .A(n10858), .Y(n5440) );
  CLKBUFX2TS U11844 ( .A(n9744), .Y(n1711) );
  CLKINVX1TS U11845 ( .A(n7526), .Y(n10054) );
  INVX2TS U11846 ( .A(n5478), .Y(n11263) );
  CLKBUFX2TS U11847 ( .A(n12411), .Y(n3644) );
  INVX2TS U11848 ( .A(n7186), .Y(n11059) );
  OR2X2TS U11849 ( .A(n9496), .B(n8665), .Y(n7390) );
  CLKINVX2TS U11850 ( .A(n3789), .Y(n11291) );
  AND2X2TS U11851 ( .A(n6724), .B(n6702), .Y(n5622) );
  INVX2TS U11852 ( .A(n2020), .Y(n12332) );
  INVX2TS U11853 ( .A(n7144), .Y(n12100) );
  CLKBUFX2TS U11854 ( .A(n11221), .Y(n5900) );
  INVX2TS U11855 ( .A(n10571), .Y(n10170) );
  INVX1TS U11856 ( .A(n6039), .Y(n10563) );
  CLKINVX2TS U11857 ( .A(n3692), .Y(n12405) );
  INVX2TS U11858 ( .A(n10959), .Y(n10142) );
  INVX2TS U11859 ( .A(n11117), .Y(n11572) );
  CLKINVX2TS U11860 ( .A(n11683), .Y(n9356) );
  INVX1TS U11861 ( .A(n5913), .Y(n10537) );
  INVX1TS U11862 ( .A(n7695), .Y(n11146) );
  INVX2TS U11863 ( .A(n7073), .Y(n11433) );
  CLKBUFX2TS U11864 ( .A(n12008), .Y(n3693) );
  AND2X2TS U11865 ( .A(n5103), .B(n4840), .Y(n4296) );
  INVX2TS U11866 ( .A(n10683), .Y(n11076) );
  INVX2TS U11867 ( .A(n7253), .Y(n10021) );
  INVX2TS U11868 ( .A(n4501), .Y(n10814) );
  INVX2TS U11869 ( .A(n7331), .Y(n11862) );
  CLKBUFX2TS U11870 ( .A(n10528), .Y(n1712) );
  INVX2TS U11871 ( .A(n9927), .Y(n10179) );
  CLKBUFX2TS U11872 ( .A(n10556), .Y(n1750) );
  INVX2TS U11873 ( .A(n7166), .Y(n11049) );
  INVX2TS U11874 ( .A(n10718), .Y(n11125) );
  INVX2TS U11875 ( .A(n10960), .Y(n11542) );
  CLKINVX2TS U11876 ( .A(n3667), .Y(n12538) );
  CLKBUFX2TS U11877 ( .A(n11837), .Y(n7422) );
  CLKINVX1TS U11878 ( .A(n3723), .Y(n11340) );
  CLKINVX2TS U11879 ( .A(n7077), .Y(n11777) );
  CLKINVX1TS U11880 ( .A(n7144), .Y(n12101) );
  INVX2TS U11881 ( .A(n7166), .Y(n11048) );
  INVX1TS U11882 ( .A(n5493), .Y(n12510) );
  CLKINVX2TS U11883 ( .A(n4321), .Y(n12490) );
  INVX2TS U11884 ( .A(n10957), .Y(n10141) );
  INVX2TS U11885 ( .A(n5913), .Y(n10535) );
  INVX2TS U11886 ( .A(n10566), .Y(n10162) );
  NOR2X1TS U11887 ( .A(n10401), .B(n12018), .Y(n4578) );
  INVX1TS U11888 ( .A(n7127), .Y(n11039) );
  INVX2TS U11889 ( .A(n7141), .Y(n11456) );
  CLKBUFX2TS U11890 ( .A(n11755), .Y(n3926) );
  INVX2TS U11891 ( .A(n2323), .Y(n9943) );
  INVX2TS U11892 ( .A(n3789), .Y(n11290) );
  INVX2TS U11893 ( .A(n10566), .Y(n10161) );
  INVX2TS U11894 ( .A(n7331), .Y(n11861) );
  INVX2TS U11895 ( .A(n9630), .Y(n9631) );
  INVX2TS U11896 ( .A(n7536), .Y(n10057) );
  CLKINVX2TS U11897 ( .A(n3723), .Y(n11339) );
  INVX2TS U11898 ( .A(n5544), .Y(n11311) );
  AND2X2TS U11899 ( .A(n4840), .B(n5106), .Y(n3930) );
  INVX1TS U11900 ( .A(n12577), .Y(n9638) );
  INVX1TS U11901 ( .A(n7238), .Y(n10623) );
  CLKBUFX2TS U11902 ( .A(n10271), .Y(n2358) );
  CLKBUFX2TS U11903 ( .A(n11404), .Y(n4044) );
  CLKBUFX2TS U11904 ( .A(n11761), .Y(n3662) );
  CLKINVX2TS U11905 ( .A(n7767), .Y(n11933) );
  INVX2TS U11906 ( .A(n7662), .Y(n12487) );
  CLKBUFX2TS U11907 ( .A(n10496), .Y(n5782) );
  INVX2TS U11908 ( .A(n1822), .Y(n11911) );
  CLKBUFX2TS U11909 ( .A(n11774), .Y(n3950) );
  INVX2TS U11910 ( .A(n7536), .Y(n10058) );
  INVX1TS U11911 ( .A(n10682), .Y(n11077) );
  INVX1TS U11912 ( .A(n5493), .Y(n12512) );
  INVX2TS U11913 ( .A(n1669), .Y(n11954) );
  INVX2TS U11914 ( .A(n4321), .Y(n12492) );
  CLKBUFX2TS U11915 ( .A(n11326), .Y(n3531) );
  INVX2TS U11916 ( .A(n10571), .Y(n10169) );
  INVX1TS U11917 ( .A(n5544), .Y(n11313) );
  INVX2TS U11918 ( .A(n7462), .Y(n11118) );
  INVX1TS U11919 ( .A(n3569), .Y(n10477) );
  INVX1TS U11920 ( .A(n7989), .Y(n10739) );
  INVX2TS U11921 ( .A(n12013), .Y(n9977) );
  INVX2TS U11922 ( .A(n9878), .Y(n11493) );
  AOI22X1TS U11923 ( .A0(n11693), .A1(n11234), .B0(n11209), .B1(n12504), .Y(
        n5849) );
  INVX1TS U11924 ( .A(n5580), .Y(n12535) );
  INVX2TS U11925 ( .A(n7992), .Y(n10352) );
  CLKBUFX2TS U11926 ( .A(n12170), .Y(n8231) );
  INVX1TS U11927 ( .A(n7298), .Y(n10643) );
  INVX1TS U11928 ( .A(n9877), .Y(n11492) );
  INVX1TS U11929 ( .A(n5478), .Y(n11265) );
  INVX2TS U11930 ( .A(n10975), .Y(n12054) );
  CLKINVX1TS U11931 ( .A(n9528), .Y(n12473) );
  AOI22X1TS U11932 ( .A0(n12252), .A1(n3555), .B0(n12057), .B1(n11405), .Y(
        n3545) );
  CLKBUFX2TS U11933 ( .A(n10085), .Y(n7299) );
  AOI22X1TS U11934 ( .A0(n12234), .A1(n5353), .B0(n11973), .B1(n11210), .Y(
        n5343) );
  INVX2TS U11935 ( .A(n5743), .Y(n11741) );
  INVX1TS U11936 ( .A(n7974), .Y(n11172) );
  CLKBUFX2TS U11937 ( .A(n11260), .Y(n3540) );
  INVX1TS U11938 ( .A(n3789), .Y(n11292) );
  AOI22X1TS U11939 ( .A0(n12228), .A1(n3594), .B0(n12051), .B1(n11394), .Y(
        n3584) );
  INVX2TS U11940 ( .A(n1756), .Y(n10658) );
  AOI22X1TS U11941 ( .A0(n12257), .A1(n5392), .B0(n11970), .B1(n11222), .Y(
        n5382) );
  CLKINVX2TS U11942 ( .A(n5513), .Y(n12426) );
  INVX1TS U11943 ( .A(n5367), .Y(n10441) );
  CLKBUFX2TS U11944 ( .A(n9833), .Y(n7292) );
  CLKINVX2TS U11945 ( .A(n7625), .Y(n10696) );
  INVX2TS U11946 ( .A(n7974), .Y(n11170) );
  INVX2TS U11947 ( .A(n9877), .Y(n11491) );
  CLKBUFX2TS U11948 ( .A(n10173), .Y(n5577) );
  INVX2TS U11949 ( .A(n9527), .Y(n12472) );
  INVX2TS U11950 ( .A(n7625), .Y(n10697) );
  INVX2TS U11951 ( .A(n12158), .Y(n10333) );
  INVX2TS U11952 ( .A(n7298), .Y(n10642) );
  INVX1TS U11953 ( .A(n7989), .Y(n10740) );
  INVX2TS U11954 ( .A(n12158), .Y(n10332) );
  AND2X2TS U11955 ( .A(n6639), .B(n6906), .Y(n5750) );
  CLKBUFX2TS U11956 ( .A(n11359), .Y(n5338) );
  INVX1TS U11957 ( .A(n5580), .Y(n12536) );
  AOI22X1TS U11958 ( .A0(n11461), .A1(n7215), .B0(n11784), .B1(n7066), .Y(
        n8633) );
  INVX2TS U11959 ( .A(n12011), .Y(n9978) );
  INVX2TS U11960 ( .A(n7186), .Y(n11060) );
  INVX2TS U11961 ( .A(n5580), .Y(n12537) );
  AOI22X1TS U11962 ( .A0(n12447), .A1(n9997), .B0(n10952), .B1(n11676), .Y(
        n6704) );
  AOI22X1TS U11963 ( .A0(n11678), .A1(n12575), .B0(n11696), .B1(n10835), .Y(
        n6734) );
  INVX2TS U11964 ( .A(n11027), .Y(n11604) );
  NOR2X1TS U11965 ( .A(n12375), .B(n10881), .Y(n3613) );
  INVX1TS U11966 ( .A(n12242), .Y(n9368) );
  AOI32XLTS U11967 ( .A0(n10748), .A1(n12043), .A2(n4000), .B0(n12071), .B1(
        n12377), .Y(n3998) );
  CLKINVX2TS U11968 ( .A(n3692), .Y(n12406) );
  OAI31X1TS U11969 ( .A0(n11418), .A1(n11798), .A2(n11793), .B0(n10928), .Y(
        n3509) );
  INVX1TS U11970 ( .A(n3530), .Y(n10495) );
  NOR2X1TS U11971 ( .A(n12447), .B(n11227), .Y(n5411) );
  AOI22X1TS U11972 ( .A0(n12375), .A1(n10129), .B0(n10801), .B1(n11787), .Y(
        n4905) );
  INVX2TS U11973 ( .A(n5657), .Y(n9974) );
  AOI22X1TS U11974 ( .A0(n11792), .A1(n12593), .B0(n12071), .B1(n10933), .Y(
        n4935) );
  INVX1TS U11975 ( .A(n4203), .Y(n9162) );
  CLKINVX2TS U11976 ( .A(n1810), .Y(n11590) );
  AOI22X1TS U11977 ( .A0(n11720), .A1(n11321), .B0(n11392), .B1(n12508), .Y(
        n4105) );
  CLKINVX2TS U11978 ( .A(n5447), .Y(n12418) );
  INVX1TS U11979 ( .A(n2220), .Y(n10583) );
  INVX1TS U11980 ( .A(n5328), .Y(n10423) );
  INVX2TS U11981 ( .A(n5745), .Y(n9727) );
  INVX2TS U11982 ( .A(n12082), .Y(n10026) );
  INVX1TS U11983 ( .A(n1822), .Y(n11913) );
  INVX1TS U11984 ( .A(n5984), .Y(n10545) );
  INVX2TS U11985 ( .A(n5585), .Y(n10946) );
  INVX1TS U11986 ( .A(n3643), .Y(n12031) );
  INVX1TS U11987 ( .A(n5984), .Y(n10546) );
  CLKINVX2TS U11988 ( .A(n3956), .Y(n11714) );
  INVX1TS U11989 ( .A(n10974), .Y(n12055) );
  CLKINVX2TS U11990 ( .A(n5745), .Y(n9726) );
  INVX2TS U11991 ( .A(n7767), .Y(n11934) );
  INVX1TS U11992 ( .A(n5743), .Y(n11742) );
  INVX2TS U11993 ( .A(n5580), .Y(n12534) );
  INVX2TS U11994 ( .A(n3667), .Y(n12540) );
  CLKINVX2TS U11995 ( .A(n1810), .Y(n11589) );
  INVX2TS U11996 ( .A(n9928), .Y(n10180) );
  INVX1TS U11997 ( .A(n2020), .Y(n12331) );
  INVX1TS U11998 ( .A(n2220), .Y(n10584) );
  INVX2TS U11999 ( .A(n5657), .Y(n9973) );
  INVX1TS U12000 ( .A(n5585), .Y(n10947) );
  INVX1TS U12001 ( .A(n7668), .Y(n11599) );
  INVX1TS U12002 ( .A(n10976), .Y(n12056) );
  CLKBUFX2TS U12003 ( .A(n10061), .Y(n7473) );
  CLKINVX1TS U12004 ( .A(n7974), .Y(n11171) );
  CLKINVX1TS U12005 ( .A(n11136), .Y(n11584) );
  AOI22X1TS U12006 ( .A0(n10797), .A1(n3659), .B0(n12199), .B1(n10396), .Y(
        n4843) );
  INVX2TS U12007 ( .A(n1718), .Y(n10671) );
  CLKBUFX2TS U12008 ( .A(n11365), .Y(n5377) );
  CLKBUFX2TS U12009 ( .A(n11254), .Y(n3579) );
  CLKBUFX2TS U12010 ( .A(n11950), .Y(n7281) );
  CLKBUFX2TS U12011 ( .A(n10305), .Y(n8191) );
  CLKINVX2TS U12012 ( .A(n3758), .Y(n12397) );
  CLKBUFX2TS U12013 ( .A(n9778), .Y(n6320) );
  CLKINVX2TS U12014 ( .A(n3756), .Y(n10438) );
  INVX2TS U12015 ( .A(n4203), .Y(n9161) );
  INVX2TS U12016 ( .A(n8351), .Y(n11198) );
  INVX1TS U12017 ( .A(n7486), .Y(n12634) );
  INVX1TS U12018 ( .A(n11478), .Y(n9984) );
  INVX2TS U12019 ( .A(n2150), .Y(n11537) );
  INVX1TS U12020 ( .A(n2019), .Y(n11057) );
  INVX2TS U12021 ( .A(n6167), .Y(n9375) );
  INVX2TS U12022 ( .A(n7940), .Y(n11940) );
  CLKINVX2TS U12023 ( .A(n3640), .Y(n11773) );
  CLKBUFX2TS U12024 ( .A(n11929), .Y(n2240) );
  CLKINVX2TS U12025 ( .A(n3574), .Y(n10895) );
  CLKINVX2TS U12026 ( .A(n3666), .Y(n11763) );
  INVX1TS U12027 ( .A(n2360), .Y(n10533) );
  INVX2TS U12028 ( .A(n2324), .Y(n12296) );
  INVX1TS U12029 ( .A(n1879), .Y(n12137) );
  INVX2TS U12030 ( .A(n7843), .Y(n11609) );
  INVX2TS U12031 ( .A(n3794), .Y(n11284) );
  INVX2TS U12032 ( .A(n1879), .Y(n12138) );
  INVX2TS U12033 ( .A(n7488), .Y(n11903) );
  INVX1TS U12034 ( .A(n3805), .Y(n11279) );
  INVX1TS U12035 ( .A(n2097), .Y(n9728) );
  CLKBUFX2TS U12036 ( .A(n10299), .Y(n2687) );
  INVX1TS U12037 ( .A(n1871), .Y(n11111) );
  CLKBUFX2TS U12038 ( .A(n11678), .Y(n6153) );
  INVX1TS U12039 ( .A(n5786), .Y(n12450) );
  CLKBUFX2TS U12040 ( .A(n10155), .Y(n3501) );
  INVX2TS U12041 ( .A(n5317), .Y(n12575) );
  CLKINVX2TS U12042 ( .A(n3929), .Y(n12572) );
  CLKBUFX2TS U12043 ( .A(n11893), .Y(n2380) );
  INVX2TS U12044 ( .A(n2324), .Y(n12295) );
  CLKINVX2TS U12045 ( .A(n3929), .Y(n12571) );
  CLKBUFX2TS U12046 ( .A(n10283), .Y(n1713) );
  CLKINVX2TS U12047 ( .A(n3672), .Y(n11757) );
  CLKINVX2TS U12048 ( .A(n5412), .Y(n11672) );
  CLKINVX1TS U12049 ( .A(n7685), .Y(n10713) );
  INVX2TS U12050 ( .A(n3993), .Y(n12375) );
  CLKINVX1TS U12051 ( .A(n4132), .Y(n10382) );
  CLKBUFX2TS U12052 ( .A(n11941), .Y(n2307) );
  OR2X2TS U12053 ( .A(n9448), .B(n6850), .Y(n5550) );
  INVX2TS U12054 ( .A(n5372), .Y(n10874) );
  INVX2TS U12055 ( .A(n5699), .Y(n11359) );
  INVX2TS U12056 ( .A(n5301), .Y(n10835) );
  INVX2TS U12057 ( .A(n1882), .Y(n10263) );
  CLKINVX2TS U12058 ( .A(n3649), .Y(n10866) );
  CLKBUFX2TS U12059 ( .A(n9845), .Y(n7322) );
  INVX1TS U12060 ( .A(n1863), .Y(n10272) );
  CLKBUFX2TS U12061 ( .A(n11695), .Y(n5293) );
  INVX1TS U12062 ( .A(n3596), .Y(n11394) );
  INVX2TS U12063 ( .A(n7685), .Y(n10711) );
  INVX1TS U12064 ( .A(n6167), .Y(n9376) );
  INVX2TS U12065 ( .A(n1865), .Y(n9744) );
  INVX1TS U12066 ( .A(n5786), .Y(n12448) );
  INVX2TS U12067 ( .A(n3614), .Y(n11386) );
  INVX1TS U12068 ( .A(n1879), .Y(n12139) );
  CLKINVX2TS U12069 ( .A(n10551), .Y(n11630) );
  INVX2TS U12070 ( .A(n3666), .Y(n11761) );
  INVX2TS U12071 ( .A(n1863), .Y(n10271) );
  INVX2TS U12072 ( .A(n1862), .Y(n11578) );
  CLKINVX1TS U12073 ( .A(n7334), .Y(n10660) );
  INVX2TS U12074 ( .A(n5317), .Y(n12576) );
  CLKBUFX2TS U12075 ( .A(n11515), .Y(n7495) );
  INVX2TS U12076 ( .A(n7313), .Y(n10285) );
  CLKINVX2TS U12077 ( .A(n5294), .Y(n12198) );
  INVX1TS U12078 ( .A(n3596), .Y(n11393) );
  CLKINVX2TS U12079 ( .A(n7055), .Y(n12069) );
  INVX1TS U12080 ( .A(n5630), .Y(n10497) );
  AND2X2TS U12081 ( .A(n9052), .B(n2598), .Y(n2590) );
  INVX2TS U12082 ( .A(n2535), .Y(n9700) );
  INVX2TS U12083 ( .A(n7326), .Y(n11101) );
  CLKINVX2TS U12084 ( .A(n5412), .Y(n11673) );
  CLKBUFX2TS U12085 ( .A(n11335), .Y(n5800) );
  INVX2TS U12086 ( .A(n2363), .Y(n10528) );
  INVX2TS U12087 ( .A(n7318), .Y(n11509) );
  CLKINVX2TS U12088 ( .A(n12201), .Y(n10776) );
  INVX2TS U12089 ( .A(n7648), .Y(n10061) );
  INVX2TS U12090 ( .A(n2196), .Y(n11003) );
  INVX2TS U12091 ( .A(n3835), .Y(n10429) );
  CLKBUFX2TS U12092 ( .A(n11983), .Y(n5582) );
  INVX2TS U12093 ( .A(n5412), .Y(n11671) );
  INVX2TS U12094 ( .A(n11307), .Y(n9961) );
  INVX2TS U12095 ( .A(n2013), .Y(n12554) );
  CLKINVX1TS U12096 ( .A(n3762), .Y(n10817) );
  INVX2TS U12097 ( .A(n3663), .Y(n10459) );
  INVX2TS U12098 ( .A(n5630), .Y(n10496) );
  INVX2TS U12099 ( .A(n2097), .Y(n9729) );
  CLKBUFX2TS U12100 ( .A(n10149), .Y(n6006) );
  INVX2TS U12101 ( .A(n3508), .Y(n12275) );
  INVX1TS U12102 ( .A(n1869), .Y(n12146) );
  CLKINVX1TS U12103 ( .A(n11488), .Y(n10543) );
  INVX1TS U12104 ( .A(n10385), .Y(n12066) );
  AND2X2TS U12105 ( .A(n3138), .B(n9051), .Y(n1803) );
  CLKINVX1TS U12106 ( .A(n3894), .Y(n11256) );
  INVX1TS U12107 ( .A(n5786), .Y(n12449) );
  INVX2TS U12108 ( .A(n7689), .Y(n10337) );
  OAI31X1TS U12109 ( .A0(n11208), .A1(n11684), .A2(n11679), .B0(n10841), .Y(
        n5307) );
  INVX2TS U12110 ( .A(n1838), .Y(n11899) );
  INVX2TS U12111 ( .A(n5663), .Y(n12005) );
  INVX2TS U12112 ( .A(n5317), .Y(n12574) );
  INVX2TS U12113 ( .A(n5983), .Y(n10233) );
  CLKBUFX2TS U12114 ( .A(n10342), .Y(n7655) );
  INVX2TS U12115 ( .A(n3652), .Y(n12411) );
  INVX1TS U12116 ( .A(n3805), .Y(n11280) );
  INVX2TS U12117 ( .A(n2952), .Y(n11423) );
  INVX2TS U12118 ( .A(n3803), .Y(n10805) );
  CLKINVX2TS U12119 ( .A(n10551), .Y(n11631) );
  CLKBUFX2TS U12120 ( .A(n10706), .Y(n7739) );
  INVX1TS U12121 ( .A(n5584), .Y(n10942) );
  INVX1TS U12122 ( .A(n1884), .Y(n9988) );
  CLKBUFX2TS U12123 ( .A(n10231), .Y(n1675) );
  CLKBUFX2TS U12124 ( .A(n11099), .Y(n1720) );
  INVX1TS U12125 ( .A(n5391), .Y(n12256) );
  INVX2TS U12126 ( .A(n3894), .Y(n11254) );
  CLKBUFX2TS U12127 ( .A(n10644), .Y(n2308) );
  CLKINVX1TS U12128 ( .A(n3574), .Y(n10893) );
  INVX2TS U12129 ( .A(n3803), .Y(n10804) );
  INVX2TS U12130 ( .A(n5584), .Y(n10941) );
  CLKINVX1TS U12131 ( .A(n7337), .Y(n11523) );
  CLKINVX2TS U12132 ( .A(n5755), .Y(n10198) );
  CLKINVX2TS U12133 ( .A(n1838), .Y(n11900) );
  INVX2TS U12134 ( .A(n1862), .Y(n11577) );
  INVX2TS U12135 ( .A(n5581), .Y(n12545) );
  INVX2TS U12136 ( .A(n7847), .Y(n9551) );
  OR2X2TS U12137 ( .A(n4516), .B(n9682), .Y(n4480) );
  INVX2TS U12138 ( .A(n7699), .Y(n11920) );
  INVX1TS U12139 ( .A(n1865), .Y(n9745) );
  INVX2TS U12140 ( .A(n2019), .Y(n11056) );
  INVX1TS U12141 ( .A(n3835), .Y(n10430) );
  INVX2TS U12142 ( .A(n7337), .Y(n11521) );
  CLKBUFX2TS U12143 ( .A(n10137), .Y(n3648) );
  INVX2TS U12144 ( .A(n4283), .Y(n10129) );
  CLKBUFX2TS U12145 ( .A(n10559), .Y(n5314) );
  CLKINVX2TS U12146 ( .A(n7326), .Y(n11102) );
  CLKINVX2TS U12147 ( .A(n7699), .Y(n11922) );
  INVX2TS U12148 ( .A(n1884), .Y(n9987) );
  INVX2TS U12149 ( .A(n2353), .Y(n10539) );
  INVX2TS U12150 ( .A(n2360), .Y(n10532) );
  INVX1TS U12151 ( .A(n2471), .Y(n10196) );
  CLKINVX2TS U12152 ( .A(n11987), .Y(n9671) );
  INVX1TS U12153 ( .A(n3794), .Y(n11286) );
  INVX2TS U12154 ( .A(n4081), .Y(n11993) );
  CLKINVX2TS U12155 ( .A(n7461), .Y(n11891) );
  CLKINVX2TS U12156 ( .A(n5983), .Y(n10234) );
  INVX2TS U12157 ( .A(n7940), .Y(n11938) );
  INVX1TS U12158 ( .A(n3739), .Y(n11328) );
  INVX2TS U12159 ( .A(n7461), .Y(n11892) );
  INVX2TS U12160 ( .A(n5575), .Y(n10173) );
  INVX2TS U12161 ( .A(n3752), .Y(n10827) );
  INVX2TS U12162 ( .A(n7075), .Y(n11032) );
  CLKINVX2TS U12163 ( .A(n3915), .Y(n12379) );
  INVX2TS U12164 ( .A(n4363), .Y(n9179) );
  INVX1TS U12165 ( .A(n2257), .Y(n12303) );
  CLKINVX2TS U12166 ( .A(n4001), .Y(n9929) );
  INVX2TS U12167 ( .A(n5954), .Y(n10226) );
  INVX1TS U12168 ( .A(n4081), .Y(n11995) );
  CLKBUFX2TS U12169 ( .A(n11729), .Y(n5593) );
  INVX2TS U12170 ( .A(n1932), .Y(n12132) );
  INVX2TS U12171 ( .A(n2257), .Y(n12302) );
  CLKINVX2TS U12172 ( .A(n7170), .Y(n11832) );
  CLKBUFX2TS U12173 ( .A(n10259), .Y(n1751) );
  CLKINVX2TS U12174 ( .A(n3920), .Y(n9651) );
  INVX2TS U12175 ( .A(n9624), .Y(n9496) );
  INVX1TS U12176 ( .A(n3503), .Y(n10934) );
  INVX2TS U12177 ( .A(n3593), .Y(n12228) );
  INVX1TS U12178 ( .A(n2293), .Y(n10561) );
  INVX1TS U12179 ( .A(n1942), .Y(n12123) );
  INVX1TS U12180 ( .A(n5994), .Y(n10550) );
  INVX2TS U12181 ( .A(n11296), .Y(n9909) );
  OR2X2TS U12182 ( .A(n9253), .B(n9249), .Y(n4108) );
  INVX2TS U12183 ( .A(n1925), .Y(n11567) );
  INVX2TS U12184 ( .A(n3519), .Y(n12593) );
  INVX2TS U12185 ( .A(n1926), .Y(n10248) );
  INVX1TS U12186 ( .A(n1928), .Y(n9741) );
  CLKBUFX2TS U12187 ( .A(n11224), .Y(n3757) );
  CLKBUFX2TS U12188 ( .A(n11869), .Y(n2424) );
  CLKINVX2TS U12189 ( .A(n7055), .Y(n12067) );
  INVX2TS U12190 ( .A(n11164), .Y(n11504) );
  INVX2TS U12191 ( .A(n1942), .Y(n12125) );
  INVX2TS U12192 ( .A(n1925), .Y(n11566) );
  INVX1TS U12193 ( .A(n7291), .Y(n12628) );
  INVX1TS U12194 ( .A(n7418), .Y(n10042) );
  INVX2TS U12195 ( .A(n3596), .Y(n11392) );
  INVX2TS U12196 ( .A(n1926), .Y(n10247) );
  INVX2TS U12197 ( .A(n1934), .Y(n11095) );
  INVX2TS U12198 ( .A(n1947), .Y(n9975) );
  CLKBUFX2TS U12199 ( .A(n11084), .Y(n1758) );
  CLKBUFX2TS U12200 ( .A(n11878), .Y(n7163) );
  CLKBUFX2TS U12201 ( .A(n10145), .Y(n5299) );
  INVX2TS U12202 ( .A(n5590), .Y(n11990) );
  CLKINVX2TS U12203 ( .A(n3666), .Y(n11762) );
  INVX2TS U12204 ( .A(n7408), .Y(n12149) );
  INVX1TS U12205 ( .A(n10045), .Y(n11086) );
  CLKINVX1TS U12206 ( .A(n3651), .Y(n9674) );
  INVX2TS U12207 ( .A(n3737), .Y(n10833) );
  INVX2TS U12208 ( .A(n3805), .Y(n11278) );
  INVX1TS U12209 ( .A(n1932), .Y(n12131) );
  CLKBUFX2TS U12210 ( .A(n9710), .Y(n5972) );
  CLKINVX2TS U12211 ( .A(n10384), .Y(n12064) );
  CLKBUFX2TS U12212 ( .A(n10273), .Y(n7169) );
  INVX2TS U12213 ( .A(n2123), .Y(n9725) );
  INVX2TS U12214 ( .A(n3869), .Y(n11260) );
  INVX1TS U12215 ( .A(n1942), .Y(n12124) );
  OR2X2TS U12216 ( .A(n9222), .B(n9253), .Y(n3567) );
  CLKINVX1TS U12217 ( .A(n10580), .Y(n11614) );
  INVX1TS U12218 ( .A(n2123), .Y(n9724) );
  CLKINVX1TS U12219 ( .A(n5333), .Y(n10857) );
  CLKINVX2TS U12220 ( .A(n5590), .Y(n11991) );
  CLKINVX1TS U12221 ( .A(n1901), .Y(n11877) );
  INVX2TS U12222 ( .A(n1901), .Y(n11875) );
  INVX2TS U12223 ( .A(n1932), .Y(n12130) );
  CLKINVX2TS U12224 ( .A(n4076), .Y(n10393) );
  INVX2TS U12225 ( .A(n2296), .Y(n10556) );
  INVX2TS U12226 ( .A(n3574), .Y(n10894) );
  CLKINVX1TS U12227 ( .A(n3535), .Y(n10910) );
  CLKINVX2TS U12228 ( .A(n3949), .Y(n10112) );
  INVX2TS U12229 ( .A(n7055), .Y(n12068) );
  CLKINVX2TS U12230 ( .A(n10578), .Y(n11612) );
  INVX2TS U12231 ( .A(n7171), .Y(n11837) );
  INVX1TS U12232 ( .A(n4552), .Y(n9686) );
  CLKINVX2TS U12233 ( .A(n5575), .Y(n10174) );
  INVX2TS U12234 ( .A(n10578), .Y(n11613) );
  CLKBUFX2TS U12235 ( .A(n3929), .Y(n12570) );
  INVX2TS U12236 ( .A(n3557), .Y(n11405) );
  OR2X2TS U12237 ( .A(n9252), .B(n5051), .Y(n3795) );
  CLKINVX2TS U12238 ( .A(n5663), .Y(n12007) );
  INVX1TS U12239 ( .A(n3663), .Y(n10460) );
  INVX2TS U12240 ( .A(n7161), .Y(n12107) );
  CLKBUFX2TS U12241 ( .A(n10295), .Y(n2720) );
  INVX2TS U12242 ( .A(n3728), .Y(n11333) );
  INVX2TS U12243 ( .A(n10612), .Y(n10614) );
  CLKINVX2TS U12244 ( .A(n1901), .Y(n11876) );
  CLKBUFX2TS U12245 ( .A(n11621), .Y(n7182) );
  CLKINVX1TS U12246 ( .A(n3696), .Y(n10844) );
  INVX2TS U12247 ( .A(n4132), .Y(n10381) );
  AOI22X1TS U12248 ( .A0(n12366), .A1(n11495), .B0(n11841), .B1(n10636), .Y(
        n2708) );
  INVX2TS U12249 ( .A(n1945), .Y(n10239) );
  NOR2X1TS U12250 ( .A(n10274), .B(n11814), .Y(n7174) );
  INVX2TS U12251 ( .A(n2286), .Y(n10565) );
  INVX1TS U12252 ( .A(n1947), .Y(n9976) );
  INVX2TS U12253 ( .A(n1928), .Y(n9740) );
  CLKINVX2TS U12254 ( .A(n3920), .Y(n9650) );
  INVX1TS U12255 ( .A(n2257), .Y(n12301) );
  CLKINVX2TS U12256 ( .A(n7243), .Y(n12122) );
  INVX2TS U12257 ( .A(n7940), .Y(n11939) );
  CLKBUFX2TS U12258 ( .A(n11527), .Y(n7846) );
  INVX2TS U12259 ( .A(n6306), .Y(n9778) );
  INVX1TS U12260 ( .A(n7109), .Y(n12304) );
  CLKINVX1TS U12261 ( .A(n6349), .Y(n9781) );
  INVX2TS U12262 ( .A(n6337), .Y(n9402) );
  INVX2TS U12263 ( .A(n1869), .Y(n12145) );
  CLKINVX2TS U12264 ( .A(n5294), .Y(n12197) );
  INVX1TS U12265 ( .A(n2324), .Y(n12297) );
  INVX1TS U12266 ( .A(n5301), .Y(n10836) );
  INVX2TS U12267 ( .A(n5581), .Y(n12542) );
  INVX2TS U12268 ( .A(n7418), .Y(n10041) );
  INVX1TS U12269 ( .A(n5558), .Y(n10936) );
  INVX2TS U12270 ( .A(n5724), .Y(n11365) );
  INVX2TS U12271 ( .A(n5994), .Y(n10549) );
  INVX2TS U12272 ( .A(n5755), .Y(n10197) );
  INVX2TS U12273 ( .A(n2293), .Y(n10560) );
  CLKINVX2TS U12274 ( .A(n3915), .Y(n12381) );
  INVX2TS U12275 ( .A(n5394), .Y(n11222) );
  CLKINVX1TS U12276 ( .A(n7843), .Y(n11611) );
  CLKINVX2TS U12277 ( .A(n7318), .Y(n11510) );
  INVX1TS U12278 ( .A(n11382), .Y(n10401) );
  CLKBUFX2TS U12279 ( .A(n11377), .Y(n6015) );
  CLKINVX2TS U12280 ( .A(n3640), .Y(n11775) );
  CLKINVX1TS U12281 ( .A(n7408), .Y(n12150) );
  CLKINVX2TS U12282 ( .A(n3894), .Y(n11255) );
  CLKINVX1TS U12283 ( .A(n7075), .Y(n11033) );
  CLKBUFX2TS U12284 ( .A(n9802), .Y(n7076) );
  INVX2TS U12285 ( .A(n5549), .Y(n11318) );
  CLKINVX2TS U12286 ( .A(n7699), .Y(n11921) );
  CLKINVX1TS U12287 ( .A(n5590), .Y(n11989) );
  CLKINVX2TS U12288 ( .A(n7685), .Y(n10712) );
  INVX2TS U12289 ( .A(n5786), .Y(n12447) );
  INVX2TS U12290 ( .A(n3915), .Y(n12380) );
  INVX2TS U12291 ( .A(n7075), .Y(n11031) );
  INVX2TS U12292 ( .A(n11988), .Y(n9672) );
  INVX2TS U12293 ( .A(n7208), .Y(n9809) );
  CLKINVX1TS U12294 ( .A(n5876), .Y(n10530) );
  CLKINVX2TS U12295 ( .A(n7689), .Y(n10338) );
  INVX2TS U12296 ( .A(n3640), .Y(n11774) );
  INVX1TS U12297 ( .A(n5560), .Y(n11325) );
  CLKBUFX2TS U12298 ( .A(n4466), .Y(n3583) );
  CLKINVX2TS U12299 ( .A(n7171), .Y(n11838) );
  INVX2TS U12300 ( .A(n5581), .Y(n12543) );
  CLKINVX1TS U12301 ( .A(n7847), .Y(n9552) );
  INVX1TS U12302 ( .A(n11381), .Y(n10400) );
  INVX1TS U12303 ( .A(n1969), .Y(n12340) );
  INVX2TS U12304 ( .A(n3511), .Y(n11416) );
  CLKINVX2TS U12305 ( .A(n7055), .Y(n12070) );
  CLKINVX2TS U12306 ( .A(n7408), .Y(n12148) );
  CLKINVX2TS U12307 ( .A(n3650), .Y(n9678) );
  CLKINVX2TS U12308 ( .A(n3652), .Y(n12412) );
  CLKBUFX2TS U12309 ( .A(n11545), .Y(n7068) );
  CLKINVX1TS U12310 ( .A(n4081), .Y(n11994) );
  INVX2TS U12311 ( .A(n5483), .Y(n11270) );
  CLKBUFX2TS U12312 ( .A(n10229), .Y(n6296) );
  CLKBUFX2TS U12313 ( .A(n12052), .Y(n3590) );
  INVX1TS U12314 ( .A(n4132), .Y(n10383) );
  INVX1TS U12315 ( .A(n7161), .Y(n12108) );
  INVX2TS U12316 ( .A(n3762), .Y(n10815) );
  INVX2TS U12317 ( .A(n3650), .Y(n9677) );
  INVX2TS U12318 ( .A(n7170), .Y(n11831) );
  CLKINVX1TS U12319 ( .A(n5590), .Y(n11992) );
  INVX2TS U12320 ( .A(n5355), .Y(n11210) );
  CLKINVX1TS U12321 ( .A(n7976), .Y(n11178) );
  CLKINVX1TS U12322 ( .A(n3652), .Y(n12413) );
  CLKINVX2TS U12323 ( .A(n7172), .Y(n10617) );
  OR2X2TS U12324 ( .A(n9398), .B(n6317), .Y(n5579) );
  CLKINVX1TS U12325 ( .A(n11496), .Y(n10570) );
  CLKINVX2TS U12326 ( .A(n7170), .Y(n11830) );
  INVX1TS U12327 ( .A(n5492), .Y(n10909) );
  INVX2TS U12328 ( .A(n6349), .Y(n9782) );
  CLKINVX2TS U12329 ( .A(n7172), .Y(n10618) );
  CLKINVX1TS U12330 ( .A(n1838), .Y(n11901) );
  INVX2TS U12331 ( .A(n5581), .Y(n12544) );
  CLKINVX2TS U12332 ( .A(n5932), .Y(n10541) );
  NOR2X1TS U12333 ( .A(n12052), .B(n12508), .Y(n4667) );
  CLKINVX1TS U12334 ( .A(n5372), .Y(n10873) );
  INVX1TS U12335 ( .A(n1932), .Y(n12133) );
  CLKINVX2TS U12336 ( .A(n5699), .Y(n11360) );
  INVX1TS U12337 ( .A(n7161), .Y(n12109) );
  INVX1TS U12338 ( .A(n7291), .Y(n12627) );
  INVX2TS U12339 ( .A(n10612), .Y(n10613) );
  CLKINVX2TS U12340 ( .A(n7334), .Y(n10661) );
  CLKINVX2TS U12341 ( .A(n8203), .Y(n11647) );
  INVX2TS U12342 ( .A(n3575), .Y(n10468) );
  CLKINVX1TS U12343 ( .A(n5451), .Y(n10898) );
  INVX1TS U12344 ( .A(n2492), .Y(n10516) );
  INVX1TS U12345 ( .A(n2173), .Y(n12311) );
  INVX2TS U12346 ( .A(n11259), .Y(n9958) );
  CLKINVX2TS U12347 ( .A(n7242), .Y(n11850) );
  CLKBUFX2TS U12348 ( .A(n11408), .Y(n5446) );
  INVX2TS U12349 ( .A(n4283), .Y(n10130) );
  INVX2TS U12350 ( .A(n7986), .Y(n10093) );
  CLKBUFX2TS U12351 ( .A(n11833), .Y(n2483) );
  CLKINVX1TS U12352 ( .A(n3614), .Y(n11388) );
  OR2X2TS U12353 ( .A(n9441), .B(n9437), .Y(n5852) );
  CLKINVX1TS U12354 ( .A(n4025), .Y(n12009) );
  INVX1TS U12355 ( .A(n3993), .Y(n12376) );
  CLKINVX1TS U12356 ( .A(n5825), .Y(n12027) );
  INVX2TS U12357 ( .A(n3949), .Y(n10111) );
  CLKBUFX2TS U12358 ( .A(n11971), .Y(n5388) );
  CLKINVX2TS U12359 ( .A(n1992), .Y(n11064) );
  INVX2TS U12360 ( .A(n3696), .Y(n10843) );
  INVX2TS U12361 ( .A(n1934), .Y(n11094) );
  INVX2TS U12362 ( .A(n5517), .Y(n10923) );
  INVX2TS U12363 ( .A(n5441), .Y(n10885) );
  INVX2TS U12364 ( .A(n1821), .Y(n12154) );
  INVX2TS U12365 ( .A(n3737), .Y(n10831) );
  INVX1TS U12366 ( .A(n2196), .Y(n11004) );
  NOR2X1TS U12367 ( .A(n12058), .B(n12522), .Y(n4595) );
  INVX2TS U12368 ( .A(n5825), .Y(n12025) );
  INVX2TS U12369 ( .A(n12035), .Y(n9771) );
  INVX1TS U12370 ( .A(n3728), .Y(n11334) );
  INVX2TS U12371 ( .A(n3651), .Y(n9673) );
  CLKINVX2TS U12372 ( .A(n5334), .Y(n10431) );
  CLKINVX2TS U12373 ( .A(n3536), .Y(n10485) );
  INVX1TS U12374 ( .A(n5483), .Y(n11271) );
  INVX2TS U12375 ( .A(n12002), .Y(n9669) );
  INVX2TS U12376 ( .A(n4025), .Y(n12008) );
  NOR2X1TS U12377 ( .A(n11973), .B(n12502), .Y(n6395) );
  INVX2TS U12378 ( .A(n5558), .Y(n10935) );
  INVX2TS U12379 ( .A(n7242), .Y(n11849) );
  INVX2TS U12380 ( .A(n5492), .Y(n10908) );
  NOR2X1TS U12381 ( .A(n11970), .B(n12519), .Y(n6467) );
  INVX2TS U12382 ( .A(n7465), .Y(n10306) );
  INVX1TS U12383 ( .A(n7357), .Y(n11534) );
  INVX2TS U12384 ( .A(n1969), .Y(n12339) );
  INVX2TS U12385 ( .A(n7291), .Y(n12626) );
  CLKBUFX2TS U12386 ( .A(n10266), .Y(n7130) );
  INVX1TS U12387 ( .A(n5549), .Y(n11319) );
  INVX2TS U12388 ( .A(n5451), .Y(n10896) );
  CLKINVX2TS U12389 ( .A(n10384), .Y(n12065) );
  CLKINVX2TS U12390 ( .A(n5373), .Y(n10448) );
  INVX2TS U12391 ( .A(n7964), .Y(n11950) );
  INVX2TS U12392 ( .A(n12050), .Y(n9774) );
  INVX1TS U12393 ( .A(n2173), .Y(n12310) );
  CLKBUFX2TS U12394 ( .A(n11974), .Y(n5349) );
  INVX1TS U12395 ( .A(n4025), .Y(n12010) );
  CLKINVX1TS U12396 ( .A(n5825), .Y(n12026) );
  INVX2TS U12397 ( .A(n5881), .Y(n12040) );
  CLKINVX2TS U12398 ( .A(n7109), .Y(n12307) );
  INVX1TS U12399 ( .A(n3737), .Y(n10832) );
  OR2X2TS U12400 ( .A(n9244), .B(n9240), .Y(n4052) );
  CLKINVX2TS U12401 ( .A(n1975), .Y(n10236) );
  INVX2TS U12402 ( .A(n3649), .Y(n10865) );
  CLKINVX2TS U12403 ( .A(n1992), .Y(n11063) );
  CLKBUFX2TS U12404 ( .A(n11231), .Y(n3691) );
  CLKBUFX2TS U12405 ( .A(n10049), .Y(n7591) );
  CLKBUFX2TS U12406 ( .A(n6229), .Y(n5342) );
  CLKINVX1TS U12407 ( .A(n5881), .Y(n12042) );
  CLKBUFX2TS U12408 ( .A(n10684), .Y(n2022) );
  INVX1TS U12409 ( .A(n1805), .Y(n11596) );
  CLKINVX1TS U12410 ( .A(n7590), .Y(n12171) );
  INVX2TS U12411 ( .A(n11346), .Y(n9906) );
  INVX2TS U12412 ( .A(n5306), .Y(n12209) );
  INVX1TS U12413 ( .A(n7455), .Y(n9834) );
  INVX2TS U12414 ( .A(n5391), .Y(n12255) );
  INVX1TS U12415 ( .A(n1942), .Y(n12126) );
  CLKINVX2TS U12416 ( .A(n7589), .Y(n12162) );
  INVX2TS U12417 ( .A(n3557), .Y(n11404) );
  INVX2TS U12418 ( .A(n11165), .Y(n11503) );
  OR2X2TS U12419 ( .A(n9449), .B(n9445), .Y(n5908) );
  INVX2TS U12420 ( .A(n3739), .Y(n11326) );
  CLKBUFX2TS U12421 ( .A(n11513), .Y(n2039) );
  OR2X2TS U12422 ( .A(n9215), .B(n9245), .Y(n3528) );
  CLKINVX1TS U12423 ( .A(n2013), .Y(n12555) );
  CLKBUFX2TS U12424 ( .A(n11414), .Y(n5512) );
  INVX2TS U12425 ( .A(n3686), .Y(n10855) );
  CLKINVX1TS U12426 ( .A(n5699), .Y(n11361) );
  INVX1TS U12427 ( .A(n3554), .Y(n12252) );
  CLKBUFX2TS U12428 ( .A(n10375), .Y(n3516) );
  INVX2TS U12429 ( .A(n11305), .Y(n9962) );
  INVX2TS U12430 ( .A(n1992), .Y(n11062) );
  CLKINVX2TS U12431 ( .A(n7551), .Y(n12334) );
  INVX2TS U12432 ( .A(n7590), .Y(n12170) );
  CLKINVX1TS U12433 ( .A(n7969), .Y(n10086) );
  INVX1TS U12434 ( .A(n8203), .Y(n11646) );
  INVX2TS U12435 ( .A(n2150), .Y(n11536) );
  INVX2TS U12436 ( .A(n1982), .Y(n11069) );
  INVX2TS U12437 ( .A(n7969), .Y(n10085) );
  CLKINVX1TS U12438 ( .A(n5517), .Y(n10925) );
  INVX2TS U12439 ( .A(n10046), .Y(n11087) );
  CLKINVX2TS U12440 ( .A(n7964), .Y(n11951) );
  INVX1TS U12441 ( .A(n4363), .Y(n9180) );
  INVX2TS U12442 ( .A(n7551), .Y(n12335) );
  CLKINVX1TS U12443 ( .A(n3696), .Y(n10845) );
  AND2X2TS U12444 ( .A(n9684), .B(n3321), .Y(n2066) );
  CLKINVX1TS U12445 ( .A(n7551), .Y(n12337) );
  INVX2TS U12446 ( .A(n7622), .Y(n11579) );
  CLKINVX2TS U12447 ( .A(n7244), .Y(n10627) );
  INVX2TS U12448 ( .A(n8203), .Y(n11645) );
  INVX1TS U12449 ( .A(n2360), .Y(n10534) );
  INVX1TS U12450 ( .A(n3519), .Y(n12594) );
  INVX1TS U12451 ( .A(n5560), .Y(n11324) );
  INVX2TS U12452 ( .A(n2173), .Y(n12308) );
  INVX1TS U12453 ( .A(n1879), .Y(n12140) );
  INVX2TS U12454 ( .A(n2471), .Y(n10195) );
  AND2X2TS U12455 ( .A(n9060), .B(n9685), .Y(n1989) );
  INVX2TS U12456 ( .A(n7589), .Y(n12163) );
  INVX2TS U12457 ( .A(n7461), .Y(n11890) );
  INVX2TS U12458 ( .A(n2492), .Y(n10514) );
  INVX2TS U12459 ( .A(n7592), .Y(n12342) );
  CLKINVX2TS U12460 ( .A(n3869), .Y(n11262) );
  INVX1TS U12461 ( .A(n3739), .Y(n11327) );
  CLKINVX2TS U12462 ( .A(n12049), .Y(n9775) );
  OR2X2TS U12463 ( .A(n9070), .B(n9951), .Y(n1960) );
  INVX2TS U12464 ( .A(n5549), .Y(n11317) );
  INVX2TS U12465 ( .A(n1871), .Y(n11110) );
  INVX1TS U12466 ( .A(n3993), .Y(n12377) );
  INVX1TS U12467 ( .A(n7622), .Y(n11581) );
  INVX2TS U12468 ( .A(n3519), .Y(n12592) );
  INVX2TS U12469 ( .A(n11166), .Y(n11505) );
  INVX2TS U12470 ( .A(n3503), .Y(n10933) );
  INVX1TS U12471 ( .A(n7590), .Y(n12172) );
  INVX2TS U12472 ( .A(n9090), .Y(n9091) );
  INVX1TS U12473 ( .A(n1982), .Y(n11068) );
  INVX1TS U12474 ( .A(n7589), .Y(n12165) );
  INVX2TS U12475 ( .A(n4001), .Y(n9930) );
  INVX2TS U12476 ( .A(n2638), .Y(n11816) );
  OR2X2TS U12477 ( .A(n9071), .B(n3325), .Y(n2168) );
  INVX2TS U12478 ( .A(n11257), .Y(n9957) );
  CLKINVX1TS U12479 ( .A(n3508), .Y(n12277) );
  INVX2TS U12480 ( .A(n1975), .Y(n10235) );
  INVX2TS U12481 ( .A(n3728), .Y(n11332) );
  INVX2TS U12482 ( .A(n5352), .Y(n12232) );
  INVX2TS U12483 ( .A(n7622), .Y(n11580) );
  INVX2TS U12484 ( .A(n5333), .Y(n10858) );
  CLKINVX2TS U12485 ( .A(n7976), .Y(n11177) );
  INVX2TS U12486 ( .A(n5373), .Y(n10449) );
  OR2X2TS U12487 ( .A(n9440), .B(n6792), .Y(n5484) );
  CLKINVX2TS U12488 ( .A(n5724), .Y(n11367) );
  CLKBUFX2TS U12489 ( .A(n11446), .Y(n2069) );
  INVX2TS U12490 ( .A(n3536), .Y(n10486) );
  INVX1TS U12491 ( .A(n1821), .Y(n12153) );
  INVX2TS U12492 ( .A(n5876), .Y(n10529) );
  CLKINVX2TS U12493 ( .A(n2535), .Y(n9701) );
  INVX2TS U12494 ( .A(n7455), .Y(n9833) );
  INVX2TS U12495 ( .A(n1982), .Y(n11067) );
  INVX2TS U12496 ( .A(n2638), .Y(n11815) );
  INVX1TS U12497 ( .A(n1821), .Y(n12152) );
  OR2X2TS U12498 ( .A(n9416), .B(n9441), .Y(n5326) );
  INVX1TS U12499 ( .A(n3993), .Y(n12378) );
  CLKINVX2TS U12500 ( .A(n7242), .Y(n11848) );
  INVX2TS U12501 ( .A(n5494), .Y(n11275) );
  INVX2TS U12502 ( .A(n5558), .Y(n10937) );
  CLKBUFX2TS U12503 ( .A(n4426), .Y(n3544) );
  CLKBUFX2TS U12504 ( .A(n6269), .Y(n5381) );
  INVX2TS U12505 ( .A(n5355), .Y(n11209) );
  INVX2TS U12506 ( .A(n1972), .Y(n10629) );
  CLKBUFX2TS U12507 ( .A(n10277), .Y(n7241) );
  INVX2TS U12508 ( .A(n2056), .Y(n10228) );
  CLKBUFX2TS U12509 ( .A(n9931), .Y(n1819) );
  INVX2TS U12510 ( .A(n11344), .Y(n9905) );
  CLKBUFX2TS U12511 ( .A(n10151), .Y(n4239) );
  INVX2TS U12512 ( .A(n1663), .Y(n10015) );
  CLKBUFX2TS U12513 ( .A(n11568), .Y(n7235) );
  INVX2TS U12514 ( .A(n3554), .Y(n12251) );
  CLKBUFX2TS U12515 ( .A(n10097), .Y(n7607) );
  INVX2TS U12516 ( .A(n7109), .Y(n12305) );
  INVX1TS U12517 ( .A(n5355), .Y(n11211) );
  CLKINVX2TS U12518 ( .A(n3614), .Y(n11387) );
  INVX2TS U12519 ( .A(n7357), .Y(n11533) );
  CLKBUFX2TS U12520 ( .A(n8270), .Y(n7975) );
  CLKINVX1TS U12521 ( .A(n7551), .Y(n12336) );
  INVX2TS U12522 ( .A(n2056), .Y(n10227) );
  INVX2TS U12523 ( .A(n2173), .Y(n12309) );
  INVX1TS U12524 ( .A(n7592), .Y(n12343) );
  INVX2TS U12525 ( .A(n3535), .Y(n10911) );
  INVX1TS U12526 ( .A(n2150), .Y(n11538) );
  INVX2TS U12527 ( .A(n7120), .Y(n10005) );
  INVX2TS U12528 ( .A(n5483), .Y(n11269) );
  OR2X2TS U12529 ( .A(n9245), .B(n4993), .Y(n3729) );
  CLKBUFX2TS U12530 ( .A(n10324), .Y(n7122) );
  INVX2TS U12531 ( .A(n5507), .Y(n10913) );
  INVX2TS U12532 ( .A(n7357), .Y(n11535) );
  INVX2TS U12533 ( .A(n1805), .Y(n11595) );
  INVX2TS U12534 ( .A(n5932), .Y(n10540) );
  CLKINVX1TS U12535 ( .A(n3508), .Y(n12276) );
  INVX1TS U12536 ( .A(n1969), .Y(n12341) );
  CLKINVX1TS U12537 ( .A(n3652), .Y(n12414) );
  OR2X2TS U12538 ( .A(n9425), .B(n9449), .Y(n5365) );
  CLKBUFX2TS U12539 ( .A(n11272), .Y(n3996) );
  INVX2TS U12540 ( .A(n1821), .Y(n12151) );
  INVX2TS U12541 ( .A(n2158), .Y(n11028) );
  CLKINVX2TS U12542 ( .A(n2013), .Y(n12556) );
  INVX2TS U12543 ( .A(n4076), .Y(n10392) );
  INVX2TS U12544 ( .A(n5560), .Y(n11323) );
  CLKINVX2TS U12545 ( .A(n1972), .Y(n10631) );
  INVX2TS U12546 ( .A(n1805), .Y(n11594) );
  CLKBUFX2TS U12547 ( .A(n9720), .Y(n2032) );
  INVX1TS U12548 ( .A(n3511), .Y(n11418) );
  CLKBUFX2TS U12549 ( .A(n10310), .Y(n8193) );
  INVX2TS U12550 ( .A(n7243), .Y(n12120) );
  CLKBUFX2TS U12551 ( .A(n10168), .Y(n1693) );
  CLKBUFX2TS U12552 ( .A(n11449), .Y(n7539) );
  CLKINVX1TS U12553 ( .A(n3915), .Y(n12382) );
  INVX1TS U12554 ( .A(n5494), .Y(n11276) );
  INVX2TS U12555 ( .A(n7465), .Y(n10305) );
  INVX2TS U12556 ( .A(n7976), .Y(n11176) );
  CLKINVX2TS U12557 ( .A(n7171), .Y(n11836) );
  INVX2TS U12558 ( .A(n5334), .Y(n10432) );
  INVX2TS U12559 ( .A(n4552), .Y(n9687) );
  INVX2TS U12560 ( .A(n1969), .Y(n12338) );
  CLKBUFX2TS U12561 ( .A(n11639), .Y(n7285) );
  INVX2TS U12562 ( .A(n5394), .Y(n11221) );
  INVX1TS U12563 ( .A(n5494), .Y(n11277) );
  INVX2TS U12564 ( .A(n7824), .Y(n12369) );
  CLKINVX1TS U12565 ( .A(n1936), .Y(n11090) );
  INVX2TS U12566 ( .A(n8069), .Y(n11628) );
  CLKINVX1TS U12567 ( .A(n8202), .Y(n10098) );
  INVX2TS U12568 ( .A(n3625), .Y(n12043) );
  INVX1TS U12569 ( .A(n5354), .Y(n11975) );
  INVX2TS U12570 ( .A(n8192), .Y(n11640) );
  INVX2TS U12571 ( .A(n7545), .Y(n10324) );
  INVX2TS U12572 ( .A(n5035), .Y(n9253) );
  OR2X2TS U12573 ( .A(n4462), .B(n9141), .Y(n3569) );
  INVX2TS U12574 ( .A(n1747), .Y(n12603) );
  INVX1TS U12575 ( .A(n8135), .Y(n11633) );
  OR2X2TS U12576 ( .A(n6048), .B(n6583), .Y(n6012) );
  INVX2TS U12577 ( .A(n7516), .Y(n12559) );
  AND2X2TS U12578 ( .A(n4086), .B(n5040), .Y(n3789) );
  INVX2TS U12579 ( .A(n1744), .Y(n11929) );
  INVX1TS U12580 ( .A(n3760), .Y(n12509) );
  INVX1TS U12581 ( .A(n2021), .Y(n12326) );
  INVX1TS U12582 ( .A(n12649), .Y(n12651) );
  INVX2TS U12583 ( .A(n1746), .Y(n12365) );
  CLKBUFX2TS U12584 ( .A(n3586), .Y(n12577) );
  CLKBUFX2TS U12585 ( .A(n5384), .Y(n12588) );
  INVX2TS U12586 ( .A(n3694), .Y(n12524) );
  INVX2TS U12587 ( .A(n7949), .Y(n11622) );
  INVX2TS U12588 ( .A(n1943), .Y(n10635) );
  INVX1TS U12589 ( .A(n1745), .Y(n11132) );
  CLKINVX2TS U12590 ( .A(n7316), .Y(n10656) );
  INVX2TS U12591 ( .A(n1767), .Y(n11923) );
  INVX2TS U12592 ( .A(n7140), .Y(n11450) );
  INVX1TS U12593 ( .A(n1943), .Y(n10637) );
  OR2X2TS U12594 ( .A(n9236), .B(n5098), .Y(n4501) );
  INVX1TS U12595 ( .A(n3595), .Y(n12053) );
  INVX2TS U12596 ( .A(n1761), .Y(n10295) );
  INVX2TS U12597 ( .A(n2197), .Y(n11508) );
  INVX1TS U12598 ( .A(n12015), .Y(n12016) );
  CLKINVX2TS U12599 ( .A(n7081), .Y(n11438) );
  INVX2TS U12600 ( .A(n3753), .Y(n11320) );
  CLKINVX2TS U12601 ( .A(n7081), .Y(n11439) );
  INVX2TS U12602 ( .A(n7329), .Y(n11516) );
  INVX1TS U12603 ( .A(n2188), .Y(n11519) );
  CLKINVX1TS U12604 ( .A(n7397), .Y(n12329) );
  AND2X2TS U12605 ( .A(n5886), .B(n6839), .Y(n5544) );
  INVX2TS U12606 ( .A(n5425), .Y(n11674) );
  AND2X2TS U12607 ( .A(n8272), .B(n9536), .Y(n8351) );
  INVX2TS U12608 ( .A(n2546), .Y(n9051) );
  INVX2TS U12609 ( .A(n3760), .Y(n12506) );
  CLKBUFX2TS U12610 ( .A(n10483), .Y(n5984) );
  INVX2TS U12611 ( .A(n10781), .Y(n10782) );
  INVX2TS U12612 ( .A(n2788), .Y(n9685) );
  CLKINVX2TS U12613 ( .A(n7691), .Y(n10343) );
  CLKBUFX2TS U12614 ( .A(n11873), .Y(n7127) );
  INVX1TS U12615 ( .A(n3492), .Y(n12074) );
  INVX2TS U12616 ( .A(n3556), .Y(n12057) );
  INVX2TS U12617 ( .A(n4256), .Y(n10375) );
  CLKINVX2TS U12618 ( .A(n10781), .Y(n10783) );
  INVX2TS U12619 ( .A(n7249), .Y(n10277) );
  INVX2TS U12620 ( .A(n1667), .Y(n12192) );
  INVX1TS U12621 ( .A(n7329), .Y(n11517) );
  INVX2TS U12622 ( .A(n5449), .Y(n12505) );
  INVX2TS U12623 ( .A(n12015), .Y(n12017) );
  INVX1TS U12624 ( .A(n3492), .Y(n12072) );
  OR2X2TS U12625 ( .A(n6265), .B(n9339), .Y(n5367) );
  CLKINVX2TS U12626 ( .A(n3319), .Y(n9071) );
  CLKINVX2TS U12627 ( .A(n7650), .Y(n9846) );
  INVX2TS U12628 ( .A(n3626), .Y(n10882) );
  INVX2TS U12629 ( .A(n3595), .Y(n12052) );
  INVX2TS U12630 ( .A(n1744), .Y(n11930) );
  INVX1TS U12631 ( .A(n4326), .Y(n10798) );
  INVX2TS U12632 ( .A(n1971), .Y(n12452) );
  CLKINVX2TS U12633 ( .A(n2484), .Y(n11458) );
  INVX2TS U12634 ( .A(n2788), .Y(n9684) );
  CLKINVX2TS U12635 ( .A(n7338), .Y(n11528) );
  CLKBUFX2TS U12636 ( .A(n10409), .Y(n3756) );
  INVX2TS U12637 ( .A(n10167), .Y(n10168) );
  INVX2TS U12638 ( .A(n5762), .Y(n11752) );
  INVX2TS U12639 ( .A(n7569), .Y(n11569) );
  INVX2TS U12640 ( .A(n1767), .Y(n11925) );
  INVX2TS U12641 ( .A(n2188), .Y(n11520) );
  AND2X2TS U12642 ( .A(n4475), .B(n5092), .Y(n3667) );
  INVX2TS U12643 ( .A(n4195), .Y(n11226) );
  CLKINVX2TS U12644 ( .A(n3502), .Y(n10152) );
  INVX2TS U12645 ( .A(n1944), .Y(n11871) );
  INVX2TS U12646 ( .A(n7568), .Y(n10688) );
  INVX2TS U12647 ( .A(n5312), .Y(n10840) );
  INVX2TS U12648 ( .A(n2649), .Y(n11440) );
  INVX2TS U12649 ( .A(n1745), .Y(n11130) );
  OR2X2TS U12650 ( .A(n5110), .B(n5098), .Y(n3643) );
  OR2X2TS U12651 ( .A(n9045), .B(n9697), .Y(n1669) );
  OR2X2TS U12652 ( .A(n8364), .B(n8521), .Y(n7974) );
  INVX1TS U12653 ( .A(n1981), .Y(n12624) );
  OR2X2TS U12654 ( .A(n5044), .B(n4439), .Y(n3804) );
  AND2X2TS U12655 ( .A(n9547), .B(n9849), .Y(n7649) );
  INVX1TS U12656 ( .A(n1747), .Y(n12604) );
  INVX2TS U12657 ( .A(n7902), .Y(n10734) );
  OR2X2TS U12658 ( .A(n8454), .B(n7860), .Y(n7486) );
  AND2X2TS U12659 ( .A(n9565), .B(n8272), .Y(n7462) );
  INVX2TS U12660 ( .A(n2189), .Y(n11513) );
  CLKINVX2TS U12661 ( .A(n2563), .Y(n9932) );
  INVX2TS U12662 ( .A(n2021), .Y(n12323) );
  INVX2TS U12663 ( .A(n1981), .Y(n12622) );
  INVX2TS U12664 ( .A(n1971), .Y(n12453) );
  INVX2TS U12665 ( .A(n1682), .Y(n10684) );
  OR2X2TS U12666 ( .A(n8466), .B(n7489), .Y(n7662) );
  INVX2TS U12667 ( .A(n4514), .Y(n9682) );
  INVX2TS U12668 ( .A(n2484), .Y(n11459) );
  AND2X2TS U12669 ( .A(n4117), .B(n4697), .Y(n4113) );
  CLKINVX2TS U12670 ( .A(n1682), .Y(n10685) );
  INVX2TS U12671 ( .A(n2277), .Y(n10986) );
  INVX2TS U12672 ( .A(n3760), .Y(n12508) );
  INVX2TS U12673 ( .A(n7650), .Y(n9845) );
  INVX1TS U12674 ( .A(n3831), .Y(n11268) );
  INVX1TS U12675 ( .A(n4481), .Y(n12621) );
  CLKINVX2TS U12676 ( .A(n2065), .Y(n12316) );
  INVX1TS U12677 ( .A(n3514), .Y(n10928) );
  INVX2TS U12678 ( .A(n2641), .Y(n11446) );
  INVX2TS U12679 ( .A(n1976), .Y(n10624) );
  INVX2TS U12680 ( .A(n12649), .Y(n12650) );
  CLKBUFX2TS U12681 ( .A(n10011), .Y(n2020) );
  INVX2TS U12682 ( .A(n7316), .Y(n10655) );
  INVX2TS U12683 ( .A(n2141), .Y(n11833) );
  INVX2TS U12684 ( .A(n3626), .Y(n10881) );
  INVX2TS U12685 ( .A(n3514), .Y(n10926) );
  CLKINVX2TS U12686 ( .A(n7548), .Y(n11128) );
  INVX2TS U12687 ( .A(n7329), .Y(n11515) );
  INVX1TS U12688 ( .A(n7824), .Y(n12370) );
  INVX2TS U12689 ( .A(n2217), .Y(n9720) );
  INVX2TS U12690 ( .A(n7691), .Y(n10342) );
  CLKBUFX2TS U12691 ( .A(n11800), .Y(n7238) );
  CLKINVX2TS U12692 ( .A(n5762), .Y(n11754) );
  INVX1TS U12693 ( .A(n1667), .Y(n12194) );
  INVX2TS U12694 ( .A(n4807), .Y(n10137) );
  INVX2TS U12695 ( .A(n7234), .Y(n11082) );
  INVX2TS U12696 ( .A(n3502), .Y(n10151) );
  CLKINVX2TS U12697 ( .A(n8220), .Y(n11652) );
  INVX1TS U12698 ( .A(n4195), .Y(n11225) );
  INVX2TS U12699 ( .A(n2034), .Y(n10231) );
  AND2X2TS U12700 ( .A(n9204), .B(n4475), .Y(n4321) );
  INVX1TS U12701 ( .A(n7824), .Y(n12371) );
  INVX2TS U12702 ( .A(n3319), .Y(n9070) );
  INVX1TS U12703 ( .A(n3753), .Y(n11322) );
  INVX2TS U12704 ( .A(n1946), .Y(n11084) );
  CLKBUFX2TS U12705 ( .A(n10604), .Y(n7767) );
  INVX2TS U12706 ( .A(n2563), .Y(n9931) );
  CLKINVX1TS U12707 ( .A(n7368), .Y(n11113) );
  INVX2TS U12708 ( .A(n2021), .Y(n12324) );
  INVX2TS U12709 ( .A(n7338), .Y(n11527) );
  CLKINVX2TS U12710 ( .A(n1976), .Y(n10626) );
  INVX2TS U12711 ( .A(n5300), .Y(n10149) );
  INVX1TS U12712 ( .A(n3625), .Y(n12046) );
  INVX2TS U12713 ( .A(n2065), .Y(n12315) );
  CLKINVX2TS U12714 ( .A(n7516), .Y(n12561) );
  INVX1TS U12715 ( .A(n1667), .Y(n12195) );
  AND2X2TS U12716 ( .A(n3137), .B(n9048), .Y(n1692) );
  OR2X2TS U12717 ( .A(n9044), .B(n9055), .Y(n1822) );
  INVX2TS U12718 ( .A(n3969), .Y(n10769) );
  INVX2TS U12719 ( .A(n7140), .Y(n11449) );
  CLKINVX2TS U12720 ( .A(n7368), .Y(n11114) );
  AND2X2TS U12721 ( .A(n3138), .B(n3137), .Y(n1810) );
  INVX2TS U12722 ( .A(n1667), .Y(n12193) );
  INVX2TS U12723 ( .A(n8192), .Y(n11639) );
  INVX2TS U12724 ( .A(n1944), .Y(n11869) );
  INVX2TS U12725 ( .A(n2546), .Y(n9052) );
  INVX2TS U12726 ( .A(n7249), .Y(n10278) );
  INVX2TS U12727 ( .A(n4195), .Y(n11224) );
  INVX2TS U12728 ( .A(n7273), .Y(n12641) );
  INVX2TS U12729 ( .A(n5576), .Y(n11983) );
  OR2X2TS U12730 ( .A(n7727), .B(n8478), .Y(n7331) );
  INVX2TS U12731 ( .A(n4280), .Y(n9657) );
  CLKINVX2TS U12732 ( .A(n2141), .Y(n11834) );
  INVX1TS U12733 ( .A(n2641), .Y(n11448) );
  INVX1TS U12734 ( .A(n1971), .Y(n12454) );
  INVX2TS U12735 ( .A(n2197), .Y(n11506) );
  INVX1TS U12736 ( .A(n4518), .Y(n10395) );
  INVX2TS U12737 ( .A(n7447), .Y(n10049) );
  INVX2TS U12738 ( .A(n1971), .Y(n12451) );
  INVX1TS U12739 ( .A(n2649), .Y(n11441) );
  OR2X2TS U12740 ( .A(n8466), .B(n7860), .Y(n7695) );
  INVX2TS U12741 ( .A(n3595), .Y(n12051) );
  CLKINVX2TS U12742 ( .A(n2641), .Y(n11447) );
  INVX2TS U12743 ( .A(n1904), .Y(n10259) );
  INVX2TS U12744 ( .A(n10265), .Y(n10266) );
  INVX1TS U12745 ( .A(n3753), .Y(n11321) );
  AND3X2TS U12746 ( .A(n9853), .B(n10336), .C(n9849), .Y(n7668) );
  INVX2TS U12747 ( .A(n8202), .Y(n10097) );
  INVX2TS U12748 ( .A(n5449), .Y(n12502) );
  INVX2TS U12749 ( .A(n1706), .Y(n11941) );
  INVX2TS U12750 ( .A(n6776), .Y(n9441) );
  INVX2TS U12751 ( .A(n8135), .Y(n11634) );
  INVX2TS U12752 ( .A(n3547), .Y(n12586) );
  CLKBUFX2TS U12753 ( .A(n11845), .Y(n1718) );
  AND2X2TS U12754 ( .A(n9506), .B(n9623), .Y(n7077) );
  INVX2TS U12755 ( .A(n7086), .Y(n11782) );
  INVX2TS U12756 ( .A(n1729), .Y(n11937) );
  INVX2TS U12757 ( .A(n1729), .Y(n11936) );
  INVX2TS U12758 ( .A(n5442), .Y(n11233) );
  INVX2TS U12759 ( .A(n7403), .Y(n11545) );
  AND2X2TS U12760 ( .A(n9624), .B(n9505), .Y(n7090) );
  INVX2TS U12761 ( .A(n3831), .Y(n11267) );
  INVX1TS U12762 ( .A(n1881), .Y(n11895) );
  INVX2TS U12763 ( .A(n7162), .Y(n11461) );
  CLKINVX2TS U12764 ( .A(n6316), .Y(n9398) );
  INVX1TS U12765 ( .A(n1707), .Y(n11153) );
  INVX2TS U12766 ( .A(n5384), .Y(n12590) );
  INVX2TS U12767 ( .A(n3556), .Y(n12059) );
  INVX2TS U12768 ( .A(n6061), .Y(n11408) );
  INVX1TS U12769 ( .A(n3513), .Y(n11792) );
  CLKINVX1TS U12770 ( .A(n5576), .Y(n11984) );
  INVX2TS U12771 ( .A(n7949), .Y(n11621) );
  INVX2TS U12772 ( .A(n7568), .Y(n10686) );
  INVX1TS U12773 ( .A(n7403), .Y(n11546) );
  INVX2TS U12774 ( .A(n3493), .Y(n10156) );
  INVX2TS U12775 ( .A(n7397), .Y(n12328) );
  CLKBUFX2TS U12776 ( .A(n10405), .Y(n3690) );
  INVX2TS U12777 ( .A(n4258), .Y(n10784) );
  INVX2TS U12778 ( .A(n4151), .Y(n11232) );
  INVX1TS U12779 ( .A(n5669), .Y(n12287) );
  INVX2TS U12780 ( .A(n5661), .Y(n11729) );
  INVX1TS U12781 ( .A(n7234), .Y(n11083) );
  INVX2TS U12782 ( .A(n2344), .Y(n10971) );
  INVX1TS U12783 ( .A(n4258), .Y(n10785) );
  CLKINVX2TS U12784 ( .A(n5576), .Y(n11982) );
  OR2X2TS U12785 ( .A(n4986), .B(n4399), .Y(n3738) );
  INVX2TS U12786 ( .A(n4280), .Y(n9656) );
  INVX1TS U12787 ( .A(n1709), .Y(n12600) );
  INVX2TS U12788 ( .A(n7081), .Y(n11437) );
  AND2X2TS U12789 ( .A(n5861), .B(n6425), .Y(n5857) );
  CLKBUFX2TS U12790 ( .A(n11426), .Y(n7186) );
  INVX1TS U12791 ( .A(n3820), .Y(n10800) );
  INVX2TS U12792 ( .A(n5393), .Y(n11971) );
  INVX2TS U12793 ( .A(n3821), .Y(n11273) );
  INVX1TS U12794 ( .A(n8069), .Y(n11629) );
  INVX2TS U12795 ( .A(n5345), .Y(n12582) );
  INVX2TS U12796 ( .A(n5626), .Y(n11342) );
  CLKBUFX2TS U12797 ( .A(n10586), .Y(n5511) );
  INVX1TS U12798 ( .A(n3556), .Y(n12058) );
  CLKINVX2TS U12799 ( .A(n7338), .Y(n11529) );
  INVX1TS U12800 ( .A(n3625), .Y(n12044) );
  INVX2TS U12801 ( .A(n6105), .Y(n11415) );
  INVX2TS U12802 ( .A(n3694), .Y(n12522) );
  INVX1TS U12803 ( .A(n1708), .Y(n12374) );
  INVX1TS U12804 ( .A(n3514), .Y(n10927) );
  CLKINVX1TS U12805 ( .A(n7516), .Y(n12560) );
  INVX2TS U12806 ( .A(n7392), .Y(n11878) );
  INVX2TS U12807 ( .A(n5515), .Y(n12520) );
  INVX2TS U12808 ( .A(n1881), .Y(n11894) );
  OR2X2TS U12809 ( .A(n6843), .B(n6242), .Y(n5559) );
  INVX2TS U12810 ( .A(n5354), .Y(n11973) );
  AND2X2TS U12811 ( .A(n9523), .B(n9607), .Y(n7131) );
  INVX1TS U12812 ( .A(n3547), .Y(n12587) );
  CLKBUFX2TS U12813 ( .A(n11764), .Y(n7393) );
  OR2X2TS U12814 ( .A(n6785), .B(n6202), .Y(n5493) );
  INVX2TS U12815 ( .A(n5449), .Y(n12504) );
  INVX2TS U12816 ( .A(n5393), .Y(n11970) );
  INVX2TS U12817 ( .A(n7135), .Y(n11806) );
  INVX1TS U12818 ( .A(n2344), .Y(n10973) );
  INVX1TS U12819 ( .A(n6061), .Y(n11409) );
  INVX1TS U12820 ( .A(n5515), .Y(n12519) );
  INVX1TS U12821 ( .A(n7466), .Y(n10311) );
  INVX2TS U12822 ( .A(n6061), .Y(n11407) );
  INVX2TS U12823 ( .A(n3627), .Y(n11786) );
  CLKBUFX2TS U12824 ( .A(n10582), .Y(n5445) );
  AND2X2TS U12825 ( .A(n4061), .B(n4625), .Y(n4057) );
  INVX1TS U12826 ( .A(n1946), .Y(n11085) );
  INVX1TS U12827 ( .A(n1944), .Y(n11870) );
  CLKINVX2TS U12828 ( .A(n5661), .Y(n11730) );
  INVX2TS U12829 ( .A(n5354), .Y(n11974) );
  INVX2TS U12830 ( .A(n5423), .Y(n11668) );
  INVX2TS U12831 ( .A(n7177), .Y(n10274) );
  CLKINVX2TS U12832 ( .A(n7397), .Y(n12327) );
  INVX2TS U12833 ( .A(n1841), .Y(n10283) );
  OR2X2TS U12834 ( .A(n6351), .B(n6900), .Y(n5743) );
  CLKINVX2TS U12835 ( .A(n8220), .Y(n11653) );
  INVX2TS U12836 ( .A(n1873), .Y(n11104) );
  INVX2TS U12837 ( .A(n1709), .Y(n12599) );
  INVX1TS U12838 ( .A(n1708), .Y(n12373) );
  INVX2TS U12839 ( .A(n1723), .Y(n10299) );
  INVX1TS U12840 ( .A(n7273), .Y(n12643) );
  CLKINVX2TS U12841 ( .A(n5661), .Y(n11728) );
  INVX1TS U12842 ( .A(n7273), .Y(n12642) );
  INVX2TS U12843 ( .A(n5290), .Y(n11695) );
  INVX2TS U12844 ( .A(n5424), .Y(n11228) );
  INVX2TS U12845 ( .A(n5311), .Y(n11678) );
  INVX1TS U12846 ( .A(n5393), .Y(n11972) );
  INVX2TS U12847 ( .A(n5615), .Y(n10951) );
  INVX1TS U12848 ( .A(n3831), .Y(n11266) );
  INVX2TS U12849 ( .A(n1880), .Y(n10644) );
  INVX1TS U12850 ( .A(n5626), .Y(n11341) );
  INVX2TS U12851 ( .A(n3820), .Y(n10799) );
  INVX2TS U12852 ( .A(n1708), .Y(n12372) );
  INVX1TS U12853 ( .A(n5290), .Y(n11697) );
  INVX2TS U12854 ( .A(n4151), .Y(n11230) );
  INVX1TS U12855 ( .A(n5778), .Y(n11379) );
  INVX1TS U12856 ( .A(n5424), .Y(n11229) );
  INVX2TS U12857 ( .A(n8220), .Y(n11654) );
  INVX1TS U12858 ( .A(n1873), .Y(n11105) );
  INVX1TS U12859 ( .A(n1873), .Y(n11106) );
  INVX2TS U12860 ( .A(n5616), .Y(n11335) );
  CLKBUFX2TS U12861 ( .A(n10750), .Y(n7298) );
  INVX2TS U12862 ( .A(n1706), .Y(n11943) );
  CLKBUFX2TS U12863 ( .A(n11944), .Y(n7625) );
  INVX2TS U12864 ( .A(n6050), .Y(n9997) );
  INVX1TS U12865 ( .A(n1883), .Y(n11100) );
  INVX2TS U12866 ( .A(n3513), .Y(n11793) );
  INVX1TS U12867 ( .A(n1841), .Y(n10284) );
  INVX2TS U12868 ( .A(n1729), .Y(n11935) );
  INVX2TS U12869 ( .A(n6024), .Y(n10559) );
  INVX1TS U12870 ( .A(n5508), .Y(n11283) );
  INVX2TS U12871 ( .A(n3492), .Y(n12071) );
  INVX2TS U12872 ( .A(n6316), .Y(n9397) );
  INVX1TS U12873 ( .A(n1723), .Y(n10300) );
  INVX1TS U12874 ( .A(n1707), .Y(n11154) );
  INVX1TS U12875 ( .A(n1706), .Y(n11942) );
  INVX1TS U12876 ( .A(n4258), .Y(n10786) );
  INVX1TS U12877 ( .A(n5312), .Y(n10842) );
  INVX1TS U12878 ( .A(n2344), .Y(n10972) );
  INVX2TS U12879 ( .A(n1883), .Y(n11099) );
  INVX2TS U12880 ( .A(n6161), .Y(n9766) );
  INVX2TS U12881 ( .A(n5424), .Y(n11227) );
  INVX1TS U12882 ( .A(n3556), .Y(n12060) );
  INVX1TS U12883 ( .A(n5384), .Y(n12591) );
  INVX2TS U12884 ( .A(n1709), .Y(n12598) );
  OR2X2TS U12885 ( .A(n9226), .B(n4783), .Y(n4272) );
  INVX1TS U12886 ( .A(n3626), .Y(n10883) );
  CLKINVX2TS U12887 ( .A(n6161), .Y(n9767) );
  CLKINVX2TS U12888 ( .A(n5300), .Y(n10150) );
  INVX1TS U12889 ( .A(n5626), .Y(n11343) );
  INVX1TS U12890 ( .A(n3694), .Y(n12523) );
  INVX2TS U12891 ( .A(n6047), .Y(n9747) );
  INVX1TS U12892 ( .A(n3760), .Y(n12507) );
  OR2X2TS U12893 ( .A(n6225), .B(n9322), .Y(n5328) );
  CLKBUFX2TS U12894 ( .A(n10690), .Y(n2220) );
  CLKBUFX2TS U12895 ( .A(n10744), .Y(n7989) );
  INVX2TS U12896 ( .A(n5309), .Y(n11206) );
  INVX2TS U12897 ( .A(n2197), .Y(n11507) );
  INVX2TS U12898 ( .A(n1881), .Y(n11893) );
  INVX2TS U12899 ( .A(n6047), .Y(n9746) );
  INVX2TS U12900 ( .A(n1707), .Y(n11152) );
  INVX2TS U12901 ( .A(n6105), .Y(n11413) );
  AND2X2TS U12902 ( .A(n5830), .B(n6781), .Y(n5478) );
  INVX1TS U12903 ( .A(n2021), .Y(n12325) );
  INVX2TS U12904 ( .A(n3493), .Y(n10155) );
  INVX2TS U12905 ( .A(n5515), .Y(n12518) );
  INVX2TS U12906 ( .A(n9801), .Y(n9802) );
  INVX2TS U12907 ( .A(n5778), .Y(n11377) );
  INVX2TS U12908 ( .A(n7516), .Y(n12558) );
  CLKBUFX2TS U12909 ( .A(n11539), .Y(n7073) );
  INVX2TS U12910 ( .A(n5291), .Y(n10146) );
  INVX1TS U12911 ( .A(n1880), .Y(n10645) );
  INVX1TS U12912 ( .A(n5312), .Y(n10841) );
  INVX2TS U12913 ( .A(n1744), .Y(n11931) );
  INVX1TS U12914 ( .A(n7086), .Y(n11784) );
  CLKBUFX2TS U12915 ( .A(n3547), .Y(n12584) );
  INVX2TS U12916 ( .A(n1747), .Y(n12602) );
  INVX1TS U12917 ( .A(n8069), .Y(n11627) );
  INVX2TS U12918 ( .A(n7368), .Y(n11112) );
  CLKINVX1TS U12919 ( .A(n3969), .Y(n10770) );
  INVX1TS U12920 ( .A(n5616), .Y(n11337) );
  INVX2TS U12921 ( .A(n5669), .Y(n12285) );
  INVX2TS U12922 ( .A(n5425), .Y(n11675) );
  INVX1TS U12923 ( .A(n2277), .Y(n10987) );
  CLKBUFX2TS U12924 ( .A(n11419), .Y(n7166) );
  INVX2TS U12925 ( .A(n1746), .Y(n12366) );
  INVX2TS U12926 ( .A(n6105), .Y(n11414) );
  AND2X2TS U12927 ( .A(n8603), .B(n9524), .Y(n7144) );
  INVX2TS U12928 ( .A(n1761), .Y(n10296) );
  INVX2TS U12929 ( .A(n4481), .Y(n12620) );
  INVX2TS U12930 ( .A(n5508), .Y(n11281) );
  AND2X2TS U12931 ( .A(n4030), .B(n4982), .Y(n3723) );
  INVX1TS U12932 ( .A(n7569), .Y(n11570) );
  INVX2TS U12933 ( .A(n4326), .Y(n10796) );
  CLKINVX2TS U12934 ( .A(n3969), .Y(n10771) );
  INVX2TS U12935 ( .A(n5616), .Y(n11336) );
  INVX2TS U12936 ( .A(n7569), .Y(n11568) );
  CLKBUFX2TS U12937 ( .A(n10517), .Y(n5585) );
  INVX2TS U12938 ( .A(n5291), .Y(n10145) );
  INVX2TS U12939 ( .A(n7177), .Y(n10273) );
  INVX2TS U12940 ( .A(n7466), .Y(n10310) );
  INVX1TS U12941 ( .A(n7392), .Y(n11880) );
  INVX2TS U12942 ( .A(n4518), .Y(n10396) );
  INVX2TS U12943 ( .A(n4977), .Y(n9244) );
  INVX1TS U12944 ( .A(n5615), .Y(n10952) );
  CLKBUFX2TS U12945 ( .A(n11839), .Y(n1756) );
  INVX2TS U12946 ( .A(n6050), .Y(n9998) );
  INVX1TS U12947 ( .A(n1745), .Y(n11131) );
  INVX2TS U12948 ( .A(n1767), .Y(n11924) );
  CLKBUFX2TS U12949 ( .A(n12075), .Y(n7512) );
  INVX2TS U12950 ( .A(n3821), .Y(n11272) );
  INVX2TS U12951 ( .A(n6834), .Y(n9449) );
  INVX1TS U12952 ( .A(n2277), .Y(n10988) );
  INVX2TS U12953 ( .A(n3687), .Y(n11368) );
  INVX1TS U12954 ( .A(n1747), .Y(n12605) );
  INVX2TS U12955 ( .A(n1936), .Y(n11089) );
  OR2X2TS U12956 ( .A(n4422), .B(n9129), .Y(n3530) );
  INVX2TS U12957 ( .A(n12631), .Y(n10298) );
  INVX2TS U12958 ( .A(n1936), .Y(n11088) );
  AND2X2TS U12959 ( .A(n4475), .B(n4532), .Y(n3956) );
  OR2X2TS U12960 ( .A(n6534), .B(n6583), .Y(n6039) );
  INVX2TS U12961 ( .A(n5959), .Y(n10229) );
  CLKBUFX2TS U12962 ( .A(n10033), .Y(n7141) );
  AND2X2TS U12963 ( .A(n5917), .B(n6497), .Y(n5913) );
  INVX2TS U12964 ( .A(n4518), .Y(n10397) );
  CLKBUFX2TS U12965 ( .A(n9722), .Y(n5580) );
  INVX1TS U12966 ( .A(n5778), .Y(n11378) );
  INVX2TS U12967 ( .A(n7949), .Y(n11623) );
  CLKINVX2TS U12968 ( .A(n7447), .Y(n10050) );
  INVX2TS U12969 ( .A(n12629), .Y(n10297) );
  INVX1TS U12970 ( .A(n8135), .Y(n11635) );
  INVX2TS U12971 ( .A(n3627), .Y(n11785) );
  INVX2TS U12972 ( .A(n7392), .Y(n11879) );
  INVX2TS U12973 ( .A(n7902), .Y(n10733) );
  CLKINVX2TS U12974 ( .A(n5669), .Y(n12286) );
  INVX1TS U12975 ( .A(n5449), .Y(n12503) );
  INVX1TS U12976 ( .A(n7568), .Y(n10687) );
  INVX2TS U12977 ( .A(n4151), .Y(n11231) );
  CLKINVX2TS U12978 ( .A(n4977), .Y(n9245) );
  CLKINVX2TS U12979 ( .A(n5675), .Y(n12013) );
  INVX2TS U12980 ( .A(n6138), .Y(n10571) );
  CLKBUFX2TS U12981 ( .A(n11710), .Y(n5373) );
  OR2X2TS U12982 ( .A(n9618), .B(n8665), .Y(n7161) );
  CLKBUFX2TS U12983 ( .A(n11734), .Y(n5584) );
  INVX2TS U12984 ( .A(n1887), .Y(n11887) );
  INVX2TS U12985 ( .A(n7280), .Y(n12635) );
  INVX2TS U12986 ( .A(n1727), .Y(n11135) );
  CLKBUFX2TS U12987 ( .A(n10640), .Y(n1934) );
  INVX2TS U12988 ( .A(n3539), .Y(n12268) );
  CLKBUFX2TS U12989 ( .A(n10473), .Y(n5994) );
  INVX2TS U12990 ( .A(n6384), .Y(n10581) );
  CLKINVX1TS U12991 ( .A(n4184), .Y(n10378) );
  CLKBUFX2TS U12992 ( .A(n11574), .Y(n7622) );
  INVX1TS U12993 ( .A(n3539), .Y(n12270) );
  OR2X2TS U12994 ( .A(n9940), .B(n9068), .Y(n1862) );
  OR2X2TS U12995 ( .A(n5693), .B(n6779), .Y(n5355) );
  AND2X2TS U12996 ( .A(n9625), .B(n9561), .Y(n7170) );
  CLKINVX2TS U12997 ( .A(n1950), .Y(n11865) );
  OR2X2TS U12998 ( .A(n9053), .B(n3198), .Y(n2360) );
  OR2X2TS U12999 ( .A(n3198), .B(n9069), .Y(n1879) );
  AND2X2TS U13000 ( .A(n8545), .B(n9477), .Y(n7461) );
  CLKBUFX2TS U13001 ( .A(n11812), .Y(n7172) );
  CLKINVX1TS U13002 ( .A(n8187), .Y(n10745) );
  INVX2TS U13003 ( .A(n7079), .Y(n10599) );
  INVX2TS U13004 ( .A(n4584), .Y(n10404) );
  INVX2TS U13005 ( .A(n6094), .Y(n10566) );
  AND2X2TS U13006 ( .A(n8648), .B(n9625), .Y(n7408) );
  NOR2X1TS U13007 ( .A(n11760), .B(n10964), .Y(n6378) );
  OR2X2TS U13008 ( .A(n9053), .B(n9939), .Y(n2353) );
  OR2X2TS U13009 ( .A(n5718), .B(n6837), .Y(n5394) );
  CLKBUFX2TS U13010 ( .A(n11203), .Y(n5483) );
  INVX2TS U13011 ( .A(n5376), .Y(n12242) );
  INVX2TS U13012 ( .A(n7378), .Y(n11539) );
  INVX1TS U13013 ( .A(n8679), .Y(n9506) );
  INVX2TS U13014 ( .A(n6314), .Y(n12063) );
  CLKBUFX2TS U13015 ( .A(n10267), .Y(n2324) );
  OR2X2TS U13016 ( .A(n7404), .B(n9618), .Y(n7075) );
  INVX1TS U13017 ( .A(n1765), .Y(n11117) );
  OR2X2TS U13018 ( .A(n6785), .B(n9322), .Y(n5494) );
  AND2X2TS U13019 ( .A(n9613), .B(n10001), .Y(n7171) );
  INVX2TS U13020 ( .A(n8187), .Y(n10744) );
  OR2X2TS U13021 ( .A(n9653), .B(n9233), .Y(n3993) );
  INVX1TS U13022 ( .A(n5376), .Y(n12243) );
  INVX2TS U13023 ( .A(n7059), .Y(n11025) );
  INVX2TS U13024 ( .A(n5760), .Y(n10517) );
  INVX2TS U13025 ( .A(n7967), .Y(n9877) );
  OR2X2TS U13026 ( .A(n8602), .B(n7547), .Y(n7357) );
  OR2X2TS U13027 ( .A(n6843), .B(n9339), .Y(n5560) );
  CLKINVX2TS U13028 ( .A(n5770), .Y(n10975) );
  CLKBUFX2TS U13029 ( .A(n11410), .Y(n3728) );
  AND3X2TS U13030 ( .A(n4464), .B(n10083), .C(n4197), .Y(n3574) );
  CLKINVX1TS U13031 ( .A(n5770), .Y(n10976) );
  OR2X2TS U13032 ( .A(n4764), .B(n9652), .Y(n3519) );
  CLKBUFX2TS U13033 ( .A(n6277), .Y(n5581) );
  INVX2TS U13034 ( .A(n6384), .Y(n10582) );
  OR2X2TS U13035 ( .A(n9712), .B(n3190), .Y(n1869) );
  INVX2TS U13036 ( .A(n5633), .Y(n10957) );
  CLKINVX2TS U13037 ( .A(n5764), .Y(n12021) );
  INVX2TS U13038 ( .A(n7070), .Y(n11419) );
  CLKBUFX2TS U13039 ( .A(n11215), .Y(n5549) );
  OR2X2TS U13040 ( .A(n9742), .B(n6728), .Y(n5630) );
  AND2X2TS U13041 ( .A(n8539), .B(n9535), .Y(n7964) );
  CLKINVX1TS U13042 ( .A(n5599), .Y(n10484) );
  NOR2X1TS U13043 ( .A(n12199), .B(n11781), .Y(n4474) );
  INVX2TS U13044 ( .A(n5733), .Y(n9722) );
  INVX2TS U13045 ( .A(n1674), .Y(n10690) );
  AND2X2TS U13046 ( .A(n9623), .B(n10002), .Y(n7055) );
  AND2X2TS U13047 ( .A(n4985), .B(n9183), .Y(n4025) );
  CLKINVX2TS U13048 ( .A(n1887), .Y(n11889) );
  INVX2TS U13049 ( .A(n7072), .Y(n11426) );
  INVX2TS U13050 ( .A(n7560), .Y(n10681) );
  OR2X2TS U13051 ( .A(n9644), .B(n9241), .Y(n3737) );
  INVX2TS U13052 ( .A(n6456), .Y(n10585) );
  CLKINVX2TS U13053 ( .A(n2388), .Y(n11477) );
  CLKBUFX2TS U13054 ( .A(n10245), .Y(n5294) );
  INVX2TS U13055 ( .A(n5376), .Y(n12241) );
  CLKINVX1TS U13056 ( .A(n6094), .Y(n10568) );
  INVX1TS U13057 ( .A(n5733), .Y(n9723) );
  CLKINVX2TS U13058 ( .A(n7586), .Y(n12155) );
  CLKBUFX2TS U13059 ( .A(n11780), .Y(n3920) );
  INVX2TS U13060 ( .A(n6456), .Y(n10586) );
  CLKBUFX2TS U13061 ( .A(n11737), .Y(n3536) );
  INVX2TS U13062 ( .A(n1950), .Y(n11863) );
  INVX2TS U13063 ( .A(n7960), .Y(n11944) );
  INVX2TS U13064 ( .A(n5337), .Y(n12219) );
  OR2X2TS U13065 ( .A(n9754), .B(n9445), .Y(n5558) );
  INVX2TS U13066 ( .A(n7056), .Y(n11764) );
  INVX2TS U13067 ( .A(n5310), .Y(n11683) );
  INVX2TS U13068 ( .A(n7960), .Y(n11945) );
  OR2X2TS U13069 ( .A(n9750), .B(n9436), .Y(n5492) );
  AND2X2TS U13070 ( .A(n6784), .B(n9380), .Y(n5825) );
  INVX2TS U13071 ( .A(n7358), .Y(n10033) );
  INVX1TS U13072 ( .A(n7126), .Y(n12084) );
  INVX2TS U13073 ( .A(n7056), .Y(n11766) );
  CLKBUFX2TS U13074 ( .A(n10649), .Y(n1871) );
  INVX2TS U13075 ( .A(n3578), .Y(n12245) );
  AND2X2TS U13076 ( .A(n9477), .B(n8520), .Y(n8203) );
  INVX2TS U13077 ( .A(n4584), .Y(n10405) );
  INVX2TS U13078 ( .A(n3539), .Y(n12269) );
  CLKAND2X2TS U13079 ( .A(n6906), .B(n6905), .Y(n5590) );
  CLKAND2X2TS U13080 ( .A(n6784), .B(n6797), .Y(n5876) );
  INVX2TS U13081 ( .A(n5310), .Y(n11684) );
  OR2X2TS U13082 ( .A(n3863), .B(n4980), .Y(n3557) );
  AND2X2TS U13083 ( .A(n6842), .B(n9384), .Y(n5881) );
  INVX2TS U13084 ( .A(n5770), .Y(n10974) );
  INVX2TS U13085 ( .A(n7110), .Y(n12075) );
  INVX2TS U13086 ( .A(n4184), .Y(n10376) );
  AND3X2TS U13087 ( .A(n6227), .B(n10075), .C(n6063), .Y(n5333) );
  OR2X2TS U13088 ( .A(n8679), .B(n9617), .Y(n7940) );
  CLKINVX1TS U13089 ( .A(n7588), .Y(n9528) );
  CLKBUFX2TS U13090 ( .A(n11692), .Y(n5334) );
  INVX2TS U13091 ( .A(n2388), .Y(n11476) );
  OR2X2TS U13092 ( .A(n4986), .B(n9129), .Y(n3739) );
  AND2X2TS U13093 ( .A(n8603), .B(n9555), .Y(n7242) );
  CLKINVX1TS U13094 ( .A(n6138), .Y(n10573) );
  CLKINVX1TS U13095 ( .A(n5675), .Y(n12014) );
  OR2X2TS U13096 ( .A(n3315), .B(n9046), .Y(n2150) );
  INVX2TS U13097 ( .A(n2164), .Y(n11530) );
  INVX2TS U13098 ( .A(n4656), .Y(n10408) );
  CLKINVX2TS U13099 ( .A(n2388), .Y(n11478) );
  OR2X2TS U13100 ( .A(n3888), .B(n5038), .Y(n3596) );
  AND2X2TS U13101 ( .A(n9898), .B(n9598), .Y(n7488) );
  AND3X2TS U13102 ( .A(sa02[0]), .B(n11180), .C(n9476), .Y(n7590) );
  INVX2TS U13103 ( .A(n3954), .Y(n10781) );
  AND2X2TS U13104 ( .A(n9607), .B(n10261), .Y(n7109) );
  INVX2TS U13105 ( .A(n3512), .Y(n11798) );
  AND2X2TS U13106 ( .A(n9060), .B(n3313), .Y(n1972) );
  INVX2TS U13107 ( .A(n7113), .Y(n10604) );
  CLKINVX2TS U13108 ( .A(n7586), .Y(n12157) );
  INVX2TS U13109 ( .A(n12645), .Y(n9999) );
  CLKBUFX2TS U13110 ( .A(n12613), .Y(n1992) );
  AND3X2TS U13111 ( .A(n6267), .B(n10103), .C(n6107), .Y(n5372) );
  CLKBUFX2TS U13112 ( .A(n11398), .Y(n3794) );
  CLKINVX2TS U13113 ( .A(n2584), .Y(n9044) );
  AND2X2TS U13114 ( .A(n9546), .B(n8443), .Y(n7318) );
  CLKAND2X2TS U13115 ( .A(n8327), .B(n8479), .Y(n7685) );
  AND2X2TS U13116 ( .A(n8579), .B(n8603), .Y(n7551) );
  INVX2TS U13117 ( .A(n5675), .Y(n12011) );
  INVX2TS U13118 ( .A(n2432), .Y(n11466) );
  INVX1TS U13119 ( .A(n4228), .Y(n10372) );
  OR2X2TS U13120 ( .A(n9732), .B(n2986), .Y(n2019) );
  OR2X2TS U13121 ( .A(n9652), .B(n4929), .Y(n3835) );
  OR2X2TS U13122 ( .A(n9716), .B(n3250), .Y(n1932) );
  OR2X2TS U13123 ( .A(n9648), .B(n9248), .Y(n3803) );
  OR2X2TS U13124 ( .A(n5044), .B(n9141), .Y(n3805) );
  INVX2TS U13125 ( .A(n3578), .Y(n12244) );
  AND2X2TS U13126 ( .A(n8414), .B(n9476), .Y(n7976) );
  CLKINVX2TS U13127 ( .A(n3838), .Y(n10795) );
  INVX2TS U13128 ( .A(n2198), .Y(n11822) );
  INVX1TS U13129 ( .A(n7070), .Y(n11420) );
  INVX2TS U13130 ( .A(n2564), .Y(n9927) );
  INVX2TS U13131 ( .A(n4656), .Y(n10409) );
  OR2X2TS U13132 ( .A(n6564), .B(n9742), .Y(n5317) );
  INVX2TS U13133 ( .A(n7133), .Y(n11043) );
  OR2X2TS U13134 ( .A(n3303), .B(n9046), .Y(n2173) );
  INVX2TS U13135 ( .A(n5594), .Y(n12279) );
  INVX2TS U13136 ( .A(n5594), .Y(n12281) );
  CLKINVX2TS U13137 ( .A(n1674), .Y(n10689) );
  CLKINVX2TS U13138 ( .A(n2584), .Y(n9045) );
  INVX2TS U13139 ( .A(n7586), .Y(n12158) );
  OR2X2TS U13140 ( .A(n9055), .B(n2998), .Y(n1805) );
  OR2X2TS U13141 ( .A(n2986), .B(n3125), .Y(n1821) );
  INVX2TS U13142 ( .A(n7588), .Y(n9527) );
  CLKINVX2TS U13143 ( .A(n5633), .Y(n10959) );
  AND2X2TS U13144 ( .A(n5043), .B(n9186), .Y(n4081) );
  INVX2TS U13145 ( .A(n7321), .Y(n11856) );
  CLKINVX2TS U13146 ( .A(n12648), .Y(n10000) );
  CLKBUFX2TS U13147 ( .A(n10243), .Y(n2257) );
  OR2X2TS U13148 ( .A(n2765), .B(n9042), .Y(n2638) );
  CLKAND2X2TS U13149 ( .A(n4925), .B(n4938), .Y(n3508) );
  OR2X2TS U13150 ( .A(n11175), .B(n8491), .Y(n7291) );
  OR2X2TS U13151 ( .A(n10092), .B(n2074), .Y(n1969) );
  CLKINVX1TS U13152 ( .A(n1671), .Y(n10012) );
  OR2X2TS U13153 ( .A(n5111), .B(n9237), .Y(n3663) );
  AND3X2TS U13154 ( .A(n9593), .B(n11174), .C(n9536), .Y(n7589) );
  INVX2TS U13155 ( .A(n2480), .Y(n10960) );
  CLKINVX2TS U13156 ( .A(n7560), .Y(n10683) );
  OR2X2TS U13157 ( .A(n2557), .B(n9056), .Y(n2196) );
  INVX2TS U13158 ( .A(n1671), .Y(n10011) );
  CLKINVX1TS U13159 ( .A(n1765), .Y(n11116) );
  AND2X2TS U13160 ( .A(n9546), .B(n8470), .Y(n7326) );
  OR2X2TS U13161 ( .A(n3258), .B(n9076), .Y(n1942) );
  INVX2TS U13162 ( .A(n1765), .Y(n11115) );
  CLKBUFX2TS U13163 ( .A(n11719), .Y(n3575) );
  CLKINVX1TS U13164 ( .A(n7700), .Y(n10718) );
  AND3X2TS U13165 ( .A(n5112), .B(n9278), .C(n3947), .Y(n3652) );
  AND3X2TS U13166 ( .A(sa32[0]), .B(n10354), .C(n9049), .Y(n2013) );
  OR3X1TS U13167 ( .A(sa03[2]), .B(n9681), .C(n9952), .Y(n12649) );
  CLKINVX2TS U13168 ( .A(n8249), .Y(n10749) );
  OR2X2TS U13169 ( .A(n9043), .B(n3026), .Y(n1982) );
  INVX2TS U13170 ( .A(n6314), .Y(n12061) );
  INVX2TS U13171 ( .A(n7321), .Y(n11855) );
  INVX2TS U13172 ( .A(n5599), .Y(n10483) );
  INVX2TS U13173 ( .A(n4228), .Y(n10371) );
  INVX2TS U13174 ( .A(n3512), .Y(n11799) );
  INVX2TS U13175 ( .A(n7321), .Y(n11854) );
  INVX2TS U13176 ( .A(n8249), .Y(n10750) );
  INVX1TS U13177 ( .A(n6314), .Y(n12062) );
  OR2X2TS U13178 ( .A(n9050), .B(n9935), .Y(n2286) );
  INVX1TS U13179 ( .A(n2121), .Y(n11841) );
  INVX2TS U13180 ( .A(n7960), .Y(n11946) );
  INVX2TS U13181 ( .A(n3838), .Y(n10793) );
  CLKAND2X2TS U13182 ( .A(n5043), .B(n5056), .Y(n4132) );
  CLKINVX2TS U13183 ( .A(n7056), .Y(n11765) );
  AND3X2TS U13184 ( .A(n4424), .B(n10055), .C(n4153), .Y(n3535) );
  INVX1TS U13185 ( .A(n1950), .Y(n11864) );
  CLKINVX1TS U13186 ( .A(n7072), .Y(n11427) );
  CLKINVX1TS U13187 ( .A(n5675), .Y(n12012) );
  CLKINVX1TS U13188 ( .A(n7126), .Y(n12083) );
  INVX2TS U13189 ( .A(n5764), .Y(n12019) );
  AND2X2TS U13190 ( .A(n8574), .B(n10262), .Y(n7243) );
  OR2X2TS U13191 ( .A(n9050), .B(n3258), .Y(n2293) );
  INVX2TS U13192 ( .A(n7700), .Y(n10717) );
  INVX2TS U13193 ( .A(n5594), .Y(n12278) );
  OR2X2TS U13194 ( .A(n9935), .B(n9075), .Y(n1925) );
  OR2X2TS U13195 ( .A(n9743), .B(n9433), .Y(n5786) );
  AND2X2TS U13196 ( .A(n9597), .B(n9547), .Y(n7699) );
  INVX1TS U13197 ( .A(n5594), .Y(n12280) );
  CLKBUFX2TS U13198 ( .A(n12638), .Y(n7244) );
  INVX2TS U13199 ( .A(n7126), .Y(n12082) );
  OR2X2TS U13200 ( .A(n2661), .B(n9952), .Y(n2492) );
  CLKINVX2TS U13201 ( .A(n2164), .Y(n11531) );
  CLKBUFX2TS U13202 ( .A(n11957), .Y(n7334) );
  AND2X2TS U13203 ( .A(n9256), .B(n3947), .Y(n3649) );
  INVX2TS U13204 ( .A(n5337), .Y(n12217) );
  INVX2TS U13205 ( .A(n7124), .Y(n11800) );
  INVX2TS U13206 ( .A(n5310), .Y(n11685) );
  CLKINVX2TS U13207 ( .A(n7110), .Y(n12076) );
  INVX1TS U13208 ( .A(n7280), .Y(n12636) );
  INVX2TS U13209 ( .A(n7366), .Y(n11873) );
  CLKINVX2TS U13210 ( .A(n7079), .Y(n10600) );
  CLKINVX2TS U13211 ( .A(n7133), .Y(n11044) );
  CLKINVX2TS U13212 ( .A(n2480), .Y(n10961) );
  CLKINVX2TS U13213 ( .A(n2432), .Y(n11464) );
  INVX2TS U13214 ( .A(n9040), .Y(n10366) );
  INVX2TS U13215 ( .A(n9900), .Y(n10365) );
  INVX2TS U13216 ( .A(n8640), .Y(n9612) );
  CLKINVX2TS U13217 ( .A(n4948), .Y(n9241) );
  OR2X2TS U13218 ( .A(n9926), .B(n4922), .Y(n3627) );
  OR2X2TS U13219 ( .A(n3185), .B(n9709), .Y(n1880) );
  INVX2TS U13220 ( .A(n2540), .Y(n11452) );
  INVX2TS U13221 ( .A(n3710), .Y(n11344) );
  INVX2TS U13222 ( .A(n3075), .Y(n9059) );
  OR2X2TS U13223 ( .A(n9925), .B(n9172), .Y(n3492) );
  INVX1TS U13224 ( .A(n3499), .Y(n12548) );
  OR2X2TS U13225 ( .A(n9704), .B(n3237), .Y(n1767) );
  INVX2TS U13226 ( .A(n3635), .Y(n11780) );
  INVX1TS U13227 ( .A(n3802), .Y(n11720) );
  INVX2TS U13228 ( .A(n7694), .Y(n9546) );
  CLKINVX2TS U13229 ( .A(n2962), .Y(n9056) );
  OR2X2TS U13230 ( .A(n9698), .B(n9695), .Y(n3514) );
  OR2X2TS U13231 ( .A(n8022), .B(n8454), .Y(n7329) );
  INVX2TS U13232 ( .A(n7158), .Y(n11812) );
  INVX2TS U13233 ( .A(n7446), .Y(n10045) );
  INVX1TS U13234 ( .A(n4039), .Y(n12003) );
  INVX2TS U13235 ( .A(n8452), .Y(n9597) );
  INVX2TS U13236 ( .A(n2144), .Y(n12613) );
  INVX2TS U13237 ( .A(n6747), .Y(n9436) );
  CLKINVX2TS U13238 ( .A(n1876), .Y(n10268) );
  AND2X2TS U13239 ( .A(n9897), .B(n8470), .Y(n7338) );
  INVX2TS U13240 ( .A(n6040), .Y(n10245) );
  INVX2TS U13241 ( .A(n4948), .Y(n9240) );
  INVX2TS U13242 ( .A(n3776), .Y(n11296) );
  INVX2TS U13243 ( .A(n2748), .Y(n9046) );
  INVX2TS U13244 ( .A(n2329), .Y(n11488) );
  OR2X2TS U13245 ( .A(n3246), .B(n2848), .Y(n1944) );
  INVX2TS U13246 ( .A(n5596), .Y(n11723) );
  OR2X2TS U13247 ( .A(n9424), .B(n6268), .Y(n5515) );
  INVX2TS U13248 ( .A(n3075), .Y(n9060) );
  INVX2TS U13249 ( .A(n4246), .Y(n9652) );
  INVX2TS U13250 ( .A(n2303), .Y(n10551) );
  INVX2TS U13251 ( .A(n5673), .Y(n11734) );
  AND3X2TS U13252 ( .A(n9097), .B(n2599), .C(n2598), .Y(n1682) );
  INVX2TS U13253 ( .A(n7230), .Y(n12638) );
  CLKINVX2TS U13254 ( .A(n4734), .Y(n9226) );
  INVX2TS U13255 ( .A(n4030), .Y(n9129) );
  CLKINVX2TS U13256 ( .A(n3499), .Y(n12549) );
  OR2X2TS U13257 ( .A(n9936), .B(n9054), .Y(n1745) );
  OR2X2TS U13258 ( .A(n9789), .B(n9786), .Y(n5312) );
  INVX2TS U13259 ( .A(n5830), .Y(n9322) );
  INVX2TS U13260 ( .A(n5557), .Y(n11710) );
  INVX1TS U13261 ( .A(n4095), .Y(n11987) );
  INVX2TS U13262 ( .A(n7611), .Y(n11574) );
  INVX1TS U13263 ( .A(n7158), .Y(n11813) );
  CLKINVX2TS U13264 ( .A(n5297), .Y(n12496) );
  CLKINVX2TS U13265 ( .A(n2748), .Y(n9047) );
  INVX2TS U13266 ( .A(n5655), .Y(n10963) );
  CLKINVX2TS U13267 ( .A(n3571), .Y(n11399) );
  INVX1TS U13268 ( .A(n3635), .Y(n11779) );
  CLKINVX2TS U13269 ( .A(n2651), .Y(n9043) );
  INVX2TS U13270 ( .A(n4335), .Y(n12199) );
  CLKINVX2TS U13271 ( .A(n5673), .Y(n11736) );
  INVX1TS U13272 ( .A(n2144), .Y(n12614) );
  INVX1TS U13273 ( .A(n4095), .Y(n11988) );
  AND2X2TS U13274 ( .A(n6914), .B(n9393), .Y(n5576) );
  OR2X2TS U13275 ( .A(n3184), .B(n2924), .Y(n1709) );
  OR4X2TS U13276 ( .A(n11173), .B(n9881), .C(sa02[6]), .D(n10068), .Y(n7273)
         );
  OR2X2TS U13277 ( .A(n8664), .B(n9580), .Y(n7949) );
  INVX2TS U13278 ( .A(n8004), .Y(n11957) );
  OR2X2TS U13279 ( .A(n9940), .B(n9061), .Y(n1707) );
  OR2X2TS U13280 ( .A(n4373), .B(n4929), .Y(n4258) );
  INVX2TS U13281 ( .A(n4335), .Y(n12202) );
  OR2X2TS U13282 ( .A(n3186), .B(n2924), .Y(n1881) );
  CLKBUFX2TS U13283 ( .A(n10257), .Y(n7548) );
  INVX2TS U13284 ( .A(n8666), .Y(n9624) );
  OR2X2TS U13285 ( .A(n9699), .B(n9232), .Y(n3831) );
  AND2X2TS U13286 ( .A(n6891), .B(n9393), .Y(n5669) );
  CLKINVX2TS U13287 ( .A(n3673), .Y(n12531) );
  OR2X2TS U13288 ( .A(n9733), .B(n3128), .Y(n2197) );
  AND2X2TS U13289 ( .A(n9560), .B(n9622), .Y(n7397) );
  OR2X2TS U13290 ( .A(n7218), .B(n8664), .Y(n7403) );
  INVX2TS U13291 ( .A(n7970), .Y(n11164) );
  OR2X2TS U13292 ( .A(n9709), .B(n3177), .Y(n1729) );
  OR2X2TS U13293 ( .A(n9061), .B(n3177), .Y(n1873) );
  INVX2TS U13294 ( .A(n1987), .Y(n12097) );
  INVX2TS U13295 ( .A(n1908), .Y(n10640) );
  INVX2TS U13296 ( .A(n8452), .Y(n9598) );
  INVX1TS U13297 ( .A(n7611), .Y(n11576) );
  INVX2TS U13298 ( .A(n6805), .Y(n9444) );
  INVX2TS U13299 ( .A(n1876), .Y(n10267) );
  INVX2TS U13300 ( .A(n7727), .Y(n10077) );
  OR2X2TS U13301 ( .A(n9200), .B(n9197), .Y(n4518) );
  OR2X2TS U13302 ( .A(n8664), .B(n8628), .Y(n7086) );
  INVX1TS U13303 ( .A(n3635), .Y(n11781) );
  INVX2TS U13304 ( .A(n5895), .Y(n12050) );
  OR2X2TS U13305 ( .A(n6177), .B(n6728), .Y(n5778) );
  INVX1TS U13306 ( .A(n5557), .Y(n11712) );
  OR2X2TS U13307 ( .A(n3189), .B(n3190), .Y(n1706) );
  INVX2TS U13308 ( .A(n5465), .Y(n11257) );
  OR2X2TS U13309 ( .A(n8657), .B(n8628), .Y(n8135) );
  INVX2TS U13310 ( .A(n8599), .Y(n10261) );
  INVX2TS U13311 ( .A(n7694), .Y(n9547) );
  INVX2TS U13312 ( .A(n7988), .Y(n9566) );
  INVX2TS U13313 ( .A(n3802), .Y(n11719) );
  INVX1TS U13314 ( .A(n5895), .Y(n12048) );
  CLKINVX2TS U13315 ( .A(n7611), .Y(n11575) );
  INVX2TS U13316 ( .A(n7727), .Y(n10078) );
  INVX2TS U13317 ( .A(n8641), .Y(n9617) );
  INVX1TS U13318 ( .A(n7446), .Y(n10046) );
  INVX2TS U13319 ( .A(n7988), .Y(n9565) );
  CLKINVX2TS U13320 ( .A(n5297), .Y(n12497) );
  OR2X2TS U13321 ( .A(n9222), .B(n9649), .Y(n4195) );
  AND3X2TS U13322 ( .A(n9452), .B(n12681), .C(n5753), .Y(n5661) );
  OR2X2TS U13323 ( .A(n9695), .B(n4373), .Y(n3626) );
  AND3X2TS U13324 ( .A(n9205), .B(n11162), .C(n10309), .Y(n3969) );
  INVX2TS U13325 ( .A(n5531), .Y(n11305) );
  OR2X2TS U13326 ( .A(n3315), .B(n3026), .Y(n1971) );
  OR2X2TS U13327 ( .A(n8657), .B(n7218), .Y(n7392) );
  INVX2TS U13328 ( .A(n5886), .Y(n9339) );
  INVX1TS U13329 ( .A(n6040), .Y(n10246) );
  OR2X2TS U13330 ( .A(n9790), .B(n9432), .Y(n5626) );
  OR2X2TS U13331 ( .A(n9985), .B(n6048), .Y(n5290) );
  OR2X2TS U13332 ( .A(n3249), .B(n3250), .Y(n1744) );
  INVX1TS U13333 ( .A(n2262), .Y(n11496) );
  INVX2TS U13334 ( .A(n2651), .Y(n9042) );
  CLKINVX2TS U13335 ( .A(n7970), .Y(n11165) );
  INVX2TS U13336 ( .A(n2962), .Y(n9055) );
  OR2X2TS U13337 ( .A(n9201), .B(n5115), .Y(n4326) );
  AND2X2TS U13338 ( .A(n9067), .B(n3313), .Y(n2641) );
  CLKINVX1TS U13339 ( .A(n5369), .Y(n11217) );
  CLKINVX2TS U13340 ( .A(n3532), .Y(n11412) );
  INVX2TS U13341 ( .A(n1845), .Y(n10649) );
  INVX2TS U13342 ( .A(n2576), .Y(n9048) );
  INVX2TS U13343 ( .A(n8666), .Y(n9625) );
  INVX1TS U13344 ( .A(n5491), .Y(n11694) );
  AND2X2TS U13345 ( .A(n3316), .B(n3322), .Y(n1976) );
  INVX2TS U13346 ( .A(n2262), .Y(n11494) );
  INVX2TS U13347 ( .A(n7619), .Y(n9536) );
  AND2X2TS U13348 ( .A(n9897), .B(n8443), .Y(n7316) );
  INVX2TS U13349 ( .A(n1939), .Y(n10243) );
  AND3X2TS U13350 ( .A(n10359), .B(sa03[3]), .C(n3316), .Y(n2141) );
  INVX2TS U13351 ( .A(n6288), .Y(n11759) );
  OR2X2TS U13352 ( .A(n9786), .B(n6177), .Y(n5424) );
  INVX1TS U13353 ( .A(n5839), .Y(n12035) );
  INVX2TS U13354 ( .A(n4039), .Y(n12001) );
  OR2X2TS U13355 ( .A(n9697), .B(n2998), .Y(n1667) );
  INVX2TS U13356 ( .A(n4734), .Y(n9225) );
  OR2X2TS U13357 ( .A(n8598), .B(n8562), .Y(n7140) );
  INVX1TS U13358 ( .A(n3776), .Y(n11298) );
  INVX2TS U13359 ( .A(n4086), .Y(n9141) );
  OR2X2TS U13360 ( .A(n9233), .B(n4373), .Y(n3821) );
  OR2X2TS U13361 ( .A(n9416), .B(n9751), .Y(n6061) );
  INVX2TS U13362 ( .A(n4095), .Y(n11985) );
  OR2X2TS U13363 ( .A(n3198), .B(n9708), .Y(n1883) );
  OR2X2TS U13364 ( .A(n9842), .B(n8599), .Y(n7568) );
  OR2X2TS U13365 ( .A(n8466), .B(n8022), .Y(n7824) );
  AND2X2TS U13366 ( .A(n6911), .B(n9392), .Y(n5762) );
  CLKINVX2TS U13367 ( .A(n5465), .Y(n11258) );
  CLKINVX2TS U13368 ( .A(n5531), .Y(n11307) );
  INVX1TS U13369 ( .A(n5655), .Y(n10964) );
  OR2X2TS U13370 ( .A(n8598), .B(n9571), .Y(n7902) );
  INVX2TS U13371 ( .A(n2278), .Y(n9717) );
  INVX2TS U13372 ( .A(n4039), .Y(n12000) );
  OR2X2TS U13373 ( .A(n9986), .B(n6721), .Y(n5425) );
  OR2X2TS U13374 ( .A(n9215), .B(n9645), .Y(n4151) );
  CLKINVX1TS U13375 ( .A(n1987), .Y(n12098) );
  OR2X2TS U13376 ( .A(n9939), .B(n9708), .Y(n1708) );
  INVX1TS U13377 ( .A(n3736), .Y(n11739) );
  CLKINVX1TS U13378 ( .A(n5465), .Y(n11259) );
  OR2X2TS U13379 ( .A(n9221), .B(n4465), .Y(n3760) );
  CLKINVX2TS U13380 ( .A(n1845), .Y(n10650) );
  OR2X2TS U13381 ( .A(n9054), .B(n3237), .Y(n1936) );
  OR2X2TS U13382 ( .A(n9415), .B(n6228), .Y(n5449) );
  INVX2TS U13383 ( .A(n7619), .Y(n9535) );
  INVX1TS U13384 ( .A(n5557), .Y(n11711) );
  OR2X2TS U13385 ( .A(n8591), .B(n8562), .Y(n8069) );
  INVX2TS U13386 ( .A(n2236), .Y(n10578) );
  INVX2TS U13387 ( .A(n2345), .Y(n9713) );
  INVX2TS U13388 ( .A(n5102), .Y(n9256) );
  INVX1TS U13389 ( .A(n4399), .Y(n9183) );
  CLKINVX2TS U13390 ( .A(n1939), .Y(n10244) );
  OR2X2TS U13391 ( .A(n9645), .B(n4993), .Y(n3556) );
  INVX2TS U13392 ( .A(n5895), .Y(n12047) );
  INVX1TS U13393 ( .A(n5596), .Y(n11722) );
  INVX1TS U13394 ( .A(n4335), .Y(n12201) );
  INVX2TS U13395 ( .A(n5369), .Y(n11215) );
  INVX2TS U13396 ( .A(n2576), .Y(n9049) );
  INVX1TS U13397 ( .A(n3736), .Y(n11738) );
  AND2X2TS U13398 ( .A(n9556), .B(n9608), .Y(n7516) );
  OR2X2TS U13399 ( .A(n3245), .B(n9705), .Y(n1943) );
  INVX1TS U13400 ( .A(n2329), .Y(n11489) );
  INVX1TS U13401 ( .A(n2144), .Y(n12615) );
  CLKINVX2TS U13402 ( .A(n5330), .Y(n11204) );
  INVX2TS U13403 ( .A(n5839), .Y(n12033) );
  INVX2TS U13404 ( .A(n3532), .Y(n11410) );
  INVX2TS U13405 ( .A(n5596), .Y(n11724) );
  OR2X2TS U13406 ( .A(n9755), .B(n6850), .Y(n5393) );
  AND2X2TS U13407 ( .A(n8579), .B(n9608), .Y(n7135) );
  INVX2TS U13408 ( .A(n5330), .Y(n11203) );
  INVX2TS U13409 ( .A(n6202), .Y(n9380) );
  OR2X2TS U13410 ( .A(n9936), .B(n9705), .Y(n1746) );
  INVX2TS U13411 ( .A(n3499), .Y(n12546) );
  INVX2TS U13412 ( .A(n4039), .Y(n12002) );
  OR2X2TS U13413 ( .A(n9751), .B(n6792), .Y(n5354) );
  INVX2TS U13414 ( .A(n5297), .Y(n12494) );
  CLKINVX1TS U13415 ( .A(n3710), .Y(n11346) );
  OR2X2TS U13416 ( .A(n9433), .B(n6177), .Y(n5616) );
  OR2X2TS U13417 ( .A(n9214), .B(n4425), .Y(n3694) );
  INVX2TS U13418 ( .A(n6013), .Y(n9742) );
  INVX1TS U13419 ( .A(n6288), .Y(n11758) );
  INVX1TS U13420 ( .A(n3802), .Y(n11721) );
  INVX2TS U13421 ( .A(n5491), .Y(n11692) );
  INVX2TS U13422 ( .A(n3673), .Y(n12530) );
  INVX2TS U13423 ( .A(n3736), .Y(n11737) );
  INVX1TS U13424 ( .A(n5491), .Y(n11693) );
  INVX2TS U13425 ( .A(n2163), .Y(n9951) );
  OR2X2TS U13426 ( .A(n3258), .B(n9704), .Y(n1946) );
  OR2X2TS U13427 ( .A(n9649), .B(n5051), .Y(n3595) );
  INVX1TS U13428 ( .A(n4335), .Y(n12200) );
  AND2X2TS U13429 ( .A(n9555), .B(n8590), .Y(n7368) );
  INVX2TS U13430 ( .A(n2262), .Y(n11495) );
  CLKINVX1TS U13431 ( .A(n7970), .Y(n11166) );
  INVX2TS U13432 ( .A(n3571), .Y(n11398) );
  OR2X2TS U13433 ( .A(n9425), .B(n9755), .Y(n6105) );
  INVX2TS U13434 ( .A(n4439), .Y(n9186) );
  AND2X2TS U13435 ( .A(n8545), .B(n9893), .Y(n8192) );
  INVX1TS U13436 ( .A(n3659), .Y(n11382) );
  INVX2TS U13437 ( .A(n3659), .Y(n11381) );
  CLKINVX2TS U13438 ( .A(n6805), .Y(n9445) );
  INVX2TS U13439 ( .A(n5573), .Y(n10473) );
  OR2X2TS U13440 ( .A(n3244), .B(n2848), .Y(n1747) );
  CLKINVX1TS U13441 ( .A(n5297), .Y(n12495) );
  OR2X2TS U13442 ( .A(n8591), .B(n7369), .Y(n7569) );
  INVX1TS U13443 ( .A(n6242), .Y(n9384) );
  OR2X2TS U13444 ( .A(n2036), .B(n2998), .Y(n2021) );
  INVX1TS U13445 ( .A(n8004), .Y(n11958) );
  INVX2TS U13446 ( .A(n5006), .Y(n9248) );
  INVX2TS U13447 ( .A(n6302), .Y(n9392) );
  CLKINVX2TS U13448 ( .A(n12740), .Y(n12710) );
  CLKINVX2TS U13449 ( .A(n12734), .Y(n12728) );
  CLKINVX2TS U13450 ( .A(n12742), .Y(n12703) );
  CLKAND2X2TS U13451 ( .A(n7154), .B(n8667), .Y(n7072) );
  AND2X2TS U13452 ( .A(n6797), .B(n6775), .Y(n6094) );
  INVX2TS U13453 ( .A(n4570), .Y(n9205) );
  INVX2TS U13454 ( .A(n6063), .Y(n9751) );
  CLKINVX2TS U13455 ( .A(n10308), .Y(n9208) );
  CLKINVX2TS U13456 ( .A(n12736), .Y(n12723) );
  CLKINVX2TS U13457 ( .A(n12744), .Y(n12699) );
  CLKINVX2TS U13458 ( .A(n12742), .Y(n12704) );
  INVX2TS U13459 ( .A(n8580), .Y(n9608) );
  CLKINVX2TS U13460 ( .A(n7546), .Y(n9842) );
  CLKINVX2TS U13461 ( .A(n4765), .Y(n9699) );
  INVX2TS U13462 ( .A(n7905), .Y(n9555) );
  INVX2TS U13463 ( .A(n4546), .Y(n9200) );
  CLKINVX2TS U13464 ( .A(n6585), .Y(n9433) );
  OR2X2TS U13465 ( .A(sa22[2]), .B(n3896), .Y(n3578) );
  INVX2TS U13466 ( .A(n4545), .Y(n9196) );
  INVX2TS U13467 ( .A(n7546), .Y(n9841) );
  INVX2TS U13468 ( .A(n2429), .Y(n9935) );
  INVX2TS U13469 ( .A(n8580), .Y(n9607) );
  INVX2TS U13470 ( .A(n9816), .Y(n9429) );
  CLKINVX2TS U13471 ( .A(n12744), .Y(n12698) );
  INVX2TS U13472 ( .A(n9374), .Y(n9589) );
  INVX1TS U13473 ( .A(n7052), .Y(n12630) );
  AND2X2TS U13474 ( .A(n2086), .B(n3191), .Y(n2388) );
  AND2X2TS U13475 ( .A(n4998), .B(n4976), .Y(n4184) );
  CLKINVX2TS U13476 ( .A(n12734), .Y(n12729) );
  CLKINVX2TS U13477 ( .A(n12743), .Y(n12702) );
  INVX2TS U13478 ( .A(n4153), .Y(n9645) );
  CLKINVX2TS U13479 ( .A(n8050), .Y(n9571) );
  INVX2TS U13480 ( .A(n2410), .Y(n9061) );
  AND2X2TS U13481 ( .A(n6855), .B(n6833), .Y(n6138) );
  AND3X2TS U13482 ( .A(n9875), .B(n9871), .C(n8600), .Y(n7110) );
  OR2X2TS U13483 ( .A(n6872), .B(n6373), .Y(n6314) );
  INVX2TS U13484 ( .A(n8237), .Y(n9893) );
  OR2X2TS U13485 ( .A(n4425), .B(n4993), .Y(n4584) );
  OR2X2TS U13486 ( .A(sa12[2]), .B(n5701), .Y(n5337) );
  CLKINVX2TS U13487 ( .A(n2384), .Y(n9708) );
  CLKINVX2TS U13488 ( .A(n12739), .Y(n12712) );
  AND3X2TS U13489 ( .A(n9119), .B(n2113), .C(n3259), .Y(n1950) );
  CLKINVX2TS U13490 ( .A(n12739), .Y(n12713) );
  INVX2TS U13491 ( .A(n9538), .Y(n9420) );
  OR2X2TS U13492 ( .A(sa01[2]), .B(n5662), .Y(n5594) );
  CLKINVX2TS U13493 ( .A(n12733), .Y(n12731) );
  CLKINVX2TS U13494 ( .A(n12739), .Y(n12714) );
  INVX2TS U13495 ( .A(n9451), .Y(n9218) );
  INVX2TS U13496 ( .A(n2560), .Y(n9696) );
  OR2X2TS U13497 ( .A(n3249), .B(n3246), .Y(n1765) );
  CLKINVX2TS U13498 ( .A(n4545), .Y(n9197) );
  INVX2TS U13499 ( .A(n6302), .Y(n9393) );
  CLKINVX2TS U13500 ( .A(n12743), .Y(n12701) );
  INVX2TS U13501 ( .A(n4197), .Y(n9649) );
  AND3X2TS U13502 ( .A(n9853), .B(n10336), .C(n8443), .Y(n7700) );
  INVX2TS U13503 ( .A(n2454), .Y(n9054) );
  CLKINVX2TS U13504 ( .A(n4806), .Y(n9237) );
  CLKINVX2TS U13505 ( .A(n4546), .Y(n9201) );
  INVX2TS U13506 ( .A(n2560), .Y(n9697) );
  CLKINVX2TS U13507 ( .A(n12741), .Y(n12708) );
  CLKINVX2TS U13508 ( .A(n2428), .Y(n9704) );
  AND3X2TS U13509 ( .A(n3306), .B(n2652), .C(n2668), .Y(n2480) );
  INVX2TS U13510 ( .A(n6063), .Y(n9750) );
  AND3X2TS U13511 ( .A(n9123), .B(n2087), .C(n3199), .Y(n1887) );
  INVX1TS U13512 ( .A(n9534), .Y(n9343) );
  CLKINVX2TS U13513 ( .A(n2429), .Y(n9936) );
  INVX2TS U13514 ( .A(n6565), .Y(n9789) );
  INVX2TS U13515 ( .A(n9431), .Y(n9326) );
  CLKINVX2TS U13516 ( .A(n12741), .Y(n12707) );
  INVX2TS U13517 ( .A(n7052), .Y(n12629) );
  INVX2TS U13518 ( .A(n8649), .Y(n9622) );
  CLKINVX2TS U13519 ( .A(n12736), .Y(n12722) );
  CLKINVX2TS U13520 ( .A(n12744), .Y(n12697) );
  INVX2TS U13521 ( .A(n9370), .Y(n9585) );
  AND2X2TS U13522 ( .A(n5056), .B(n5034), .Y(n4228) );
  INVX2TS U13523 ( .A(n3100), .Y(n9063) );
  OR2X2TS U13524 ( .A(n4465), .B(n5051), .Y(n4656) );
  AND2X2TS U13525 ( .A(n2112), .B(n3251), .Y(n2432) );
  INVX2TS U13526 ( .A(n7106), .Y(n10257) );
  INVX2TS U13527 ( .A(n10732), .Y(n9593) );
  INVX2TS U13528 ( .A(n3100), .Y(n9062) );
  INVX2TS U13529 ( .A(n2384), .Y(n9709) );
  OR2X2TS U13530 ( .A(sa30[2]), .B(n5427), .Y(n5310) );
  INVX2TS U13531 ( .A(n4281), .Y(n9172) );
  INVX2TS U13532 ( .A(n9892), .Y(n9229) );
  INVX2TS U13533 ( .A(n2029), .Y(n9732) );
  INVX2TS U13534 ( .A(sa00[4]), .Y(n9193) );
  INVX2TS U13535 ( .A(n5821), .Y(n9985) );
  INVX2TS U13536 ( .A(n2428), .Y(n9705) );
  INVX2TS U13537 ( .A(n9462), .Y(n9097) );
  AND3X2TS U13538 ( .A(n9803), .B(n9799), .C(n8667), .Y(n7056) );
  INVX2TS U13539 ( .A(n4000), .Y(n9925) );
  INVX2TS U13540 ( .A(n2385), .Y(n9939) );
  INVX2TS U13541 ( .A(n4570), .Y(n9204) );
  INVX2TS U13542 ( .A(n7905), .Y(n9556) );
  OR2X2TS U13543 ( .A(n11168), .B(n3871), .Y(n3539) );
  INVX2TS U13544 ( .A(n6107), .Y(n9754) );
  INVX2TS U13545 ( .A(n8341), .Y(n9898) );
  OR2X2TS U13546 ( .A(n10350), .B(n1824), .Y(n2198) );
  OR2X2TS U13547 ( .A(n11201), .B(n5726), .Y(n5376) );
  INVX2TS U13548 ( .A(n8237), .Y(n9894) );
  OR2X2TS U13549 ( .A(n6228), .B(n6792), .Y(n6384) );
  OR2X2TS U13550 ( .A(n9892), .B(n3629), .Y(n3512) );
  CLKINVX2TS U13551 ( .A(n12741), .Y(n12706) );
  INVX2TS U13552 ( .A(n8649), .Y(n9623) );
  CLKINVX2TS U13553 ( .A(n12740), .Y(n12709) );
  INVX2TS U13554 ( .A(n9435), .Y(n9411) );
  CLKINVX2TS U13555 ( .A(n4785), .Y(n9233) );
  CLKINVX2TS U13556 ( .A(n12740), .Y(n12711) );
  INVX2TS U13557 ( .A(n4765), .Y(n9698) );
  INVX1TS U13558 ( .A(n9447), .Y(n9144) );
  INVX2TS U13559 ( .A(n7952), .Y(n9560) );
  INVX2TS U13560 ( .A(n9348), .Y(n9132) );
  CLKINVX2TS U13561 ( .A(n12733), .Y(n12730) );
  INVX2TS U13562 ( .A(n9526), .Y(n9681) );
  CLKINVX2TS U13563 ( .A(n8116), .Y(n9581) );
  INVX2TS U13564 ( .A(n3305), .Y(n9067) );
  CLKINVX2TS U13565 ( .A(n12743), .Y(n12700) );
  CLKINVX2TS U13566 ( .A(n12733), .Y(n12732) );
  CLKINVX2TS U13567 ( .A(n12736), .Y(n12721) );
  AND2X2TS U13568 ( .A(n6319), .B(n6891), .Y(n5675) );
  INVX2TS U13569 ( .A(n9345), .Y(n9452) );
  INVX2TS U13570 ( .A(n11175), .Y(n9539) );
  INVX2TS U13571 ( .A(n3305), .Y(n9066) );
  OR2X2TS U13572 ( .A(n6268), .B(n6850), .Y(n6456) );
  INVX2TS U13573 ( .A(n9351), .Y(n9211) );
  AND3X2TS U13574 ( .A(n10359), .B(sa03[3]), .C(n2167), .Y(n2164) );
  INVX2TS U13575 ( .A(n7952), .Y(n9561) );
  INVX2TS U13576 ( .A(n4153), .Y(n9644) );
  OR2X2TS U13577 ( .A(sa31[2]), .B(n7829), .Y(n7321) );
  CLKINVX2TS U13578 ( .A(n12742), .Y(n12705) );
  CLKINVX2TS U13579 ( .A(n12734), .Y(n12727) );
  INVX2TS U13580 ( .A(n8341), .Y(n9897) );
  AND3X2TS U13581 ( .A(n6911), .B(sa01[0]), .C(n10048), .Y(n5770) );
  INVX1TS U13582 ( .A(n7052), .Y(n12631) );
  AND2X2TS U13583 ( .A(n8271), .B(n8520), .Y(n8187) );
  OR2X2TS U13584 ( .A(n3189), .B(n3186), .Y(n1727) );
  AND3X2TS U13585 ( .A(sa02[0]), .B(n11180), .C(n8271), .Y(n8249) );
  INVX2TS U13586 ( .A(n4197), .Y(n9648) );
  OR2X2TS U13587 ( .A(n8523), .B(n8488), .Y(n7960) );
  CLKINVX2TS U13588 ( .A(n12745), .Y(n12696) );
  INVX2TS U13589 ( .A(n6107), .Y(n9755) );
  CLKINVX2TS U13590 ( .A(n6565), .Y(n9790) );
  INVX2TS U13591 ( .A(n11966), .Y(n11659) );
  INVX2TS U13592 ( .A(n11648), .Y(n11650) );
  INVX2TS U13593 ( .A(n9040), .Y(n11660) );
  INVX2TS U13594 ( .A(n9899), .Y(n12610) );
  INVX2TS U13595 ( .A(n9899), .Y(n12607) );
  INVX2TS U13596 ( .A(n11662), .Y(n11663) );
  INVX2TS U13597 ( .A(n11655), .Y(n11656) );
  INVX2TS U13598 ( .A(n9899), .Y(n11665) );
  INVX2TS U13599 ( .A(n9900), .Y(n12609) );
  INVX2TS U13600 ( .A(n11655), .Y(n11657) );
  INVX2TS U13601 ( .A(n11662), .Y(n11664) );
  INVX2TS U13602 ( .A(n9040), .Y(n11666) );
  INVX2TS U13603 ( .A(n9899), .Y(n10361) );
  INVX2TS U13604 ( .A(n11648), .Y(n11649) );
  CLKINVX2TS U13605 ( .A(n12735), .Y(n12724) );
  OR2X2TS U13606 ( .A(n6640), .B(n6897), .Y(n5596) );
  OR2X2TS U13607 ( .A(n3249), .B(n3244), .Y(n2262) );
  CLKINVX2TS U13608 ( .A(n12735), .Y(n12725) );
  OR2X2TS U13609 ( .A(n6872), .B(n6640), .Y(n5655) );
  INVX1TS U13610 ( .A(n12644), .Y(n12646) );
  OR2X2TS U13611 ( .A(n3189), .B(n3184), .Y(n2329) );
  INVX2TS U13612 ( .A(n12644), .Y(n12645) );
  INVX1TS U13613 ( .A(n12644), .Y(n12647) );
  AND3X2TS U13614 ( .A(n10345), .B(sa02[3]), .C(n8535), .Y(n7970) );
  AND3X2TS U13615 ( .A(n11162), .B(n10308), .C(n5092), .Y(n3659) );
  OR2X2TS U13616 ( .A(n5693), .B(n6785), .Y(n5839) );
  OR2X2TS U13617 ( .A(n3863), .B(n4986), .Y(n4039) );
  OR2X2TS U13618 ( .A(n5718), .B(n6843), .Y(n5895) );
  OR2X2TS U13619 ( .A(n3888), .B(n5044), .Y(n4095) );
  CLKINVX2TS U13620 ( .A(n12735), .Y(n12726) );
  INVX1TS U13621 ( .A(n12644), .Y(n12648) );
  OR2X2TS U13622 ( .A(n5074), .B(n5110), .Y(n4335) );
  INVX2TS U13623 ( .A(n12606), .Y(n9899) );
  CLKINVX2TS U13624 ( .A(n7991), .Y(n9882) );
  CLKINVX2TS U13625 ( .A(n8453), .Y(n9603) );
  INVX2TS U13626 ( .A(n8453), .Y(n9602) );
  INVX2TS U13627 ( .A(n7991), .Y(n9881) );
  INVX2TS U13628 ( .A(n1731), .Y(n9124) );
  INVX2TS U13629 ( .A(n7656), .Y(n9853) );
  OR4X2TS U13630 ( .A(n9792), .B(n10705), .C(sa20[7]), .D(sa20[5]), .Y(n7052)
         );
  INVX2TS U13631 ( .A(n1769), .Y(n9120) );
  OR4X2TS U13632 ( .A(sa32[7]), .B(sa32[5]), .C(n9462), .D(n10355), .Y(n12644)
         );
  INVX2TS U13633 ( .A(n10714), .Y(n10715) );
  INVX2TS U13634 ( .A(n9883), .Y(n9884) );
  INVX2TS U13635 ( .A(n9540), .Y(n9541) );
  INVX2TS U13636 ( .A(n10067), .Y(n10068) );
  INVX2TS U13637 ( .A(n10741), .Y(n10743) );
  CLKINVX2TS U13638 ( .A(n12737), .Y(n12719) );
  INVX2TS U13639 ( .A(n9823), .Y(n9824) );
  INVX2TS U13640 ( .A(n10703), .Y(n10704) );
  INVX2TS U13641 ( .A(n9847), .Y(n9848) );
  INVX2TS U13642 ( .A(n10059), .Y(n10060) );
  INVX2TS U13643 ( .A(n9887), .Y(n9888) );
  INVX2TS U13644 ( .A(n9871), .Y(n9872) );
  INVX2TS U13645 ( .A(n10099), .Y(n10100) );
  INVX2TS U13646 ( .A(n10746), .Y(n10747) );
  INVX2TS U13647 ( .A(n10075), .Y(n10076) );
  INVX2TS U13648 ( .A(n9839), .Y(n9840) );
  INVX2TS U13649 ( .A(n10079), .Y(n10080) );
  INVX2TS U13650 ( .A(n9791), .Y(n9792) );
  INVX2TS U13651 ( .A(n10071), .Y(n10072) );
  INVX1TS U13652 ( .A(n9277), .Y(n9278) );
  INVX2TS U13653 ( .A(n9787), .Y(n9788) );
  INVX2TS U13654 ( .A(n9863), .Y(n9864) );
  INVX2TS U13655 ( .A(n10103), .Y(n10104) );
  INVX2TS U13656 ( .A(n11184), .Y(n11186) );
  INVX2TS U13657 ( .A(n10307), .Y(n10308) );
  INVX2TS U13658 ( .A(n10367), .Y(n10368) );
  INVX2TS U13659 ( .A(n10051), .Y(n10052) );
  INVX2TS U13660 ( .A(n9867), .Y(n9868) );
  INVX2TS U13661 ( .A(n9799), .Y(n9800) );
  INVX2TS U13662 ( .A(n9434), .Y(n9435) );
  INVX2TS U13663 ( .A(n10055), .Y(n10056) );
  INVX2TS U13664 ( .A(n10730), .Y(n10731) );
  INVX2TS U13665 ( .A(n10083), .Y(n10084) );
  INVX2TS U13666 ( .A(n9875), .Y(n9876) );
  INVX2TS U13667 ( .A(n9815), .Y(n9816) );
  INVX2TS U13668 ( .A(n9803), .Y(n9804) );
  INVX2TS U13669 ( .A(n11189), .Y(n11191) );
  INVX2TS U13670 ( .A(n10714), .Y(n10716) );
  INVX2TS U13671 ( .A(n10322), .Y(n10323) );
  INVX2TS U13672 ( .A(n10326), .Y(n10327) );
  INVX2TS U13673 ( .A(n9430), .Y(n9431) );
  INVX2TS U13674 ( .A(n9457), .Y(n9458) );
  INVX2TS U13675 ( .A(n10312), .Y(n10314) );
  INVX2TS U13676 ( .A(n10720), .Y(n10721) );
  INVX2TS U13677 ( .A(n10035), .Y(n10036) );
  INVX2TS U13678 ( .A(n10751), .Y(n10752) );
  INVX2TS U13679 ( .A(n9544), .Y(n9545) );
  INVX2TS U13680 ( .A(n10741), .Y(n10742) );
  INVX2TS U13681 ( .A(n9831), .Y(n9832) );
  INVX2TS U13682 ( .A(n10031), .Y(n10032) );
  CLKINVX2TS U13683 ( .A(n10307), .Y(n10309) );
  INVX2TS U13684 ( .A(n9438), .Y(n9439) );
  INVX2TS U13685 ( .A(n9357), .Y(n9358) );
  INVX2TS U13686 ( .A(n11184), .Y(n11185) );
  INVX2TS U13687 ( .A(n10698), .Y(n10699) );
  INVX2TS U13688 ( .A(n10312), .Y(n10313) );
  INVX2TS U13689 ( .A(n9835), .Y(n9836) );
  CLKINVX2TS U13690 ( .A(n11173), .Y(n11174) );
  INVX2TS U13691 ( .A(n9807), .Y(n9808) );
  INVX2TS U13692 ( .A(n9891), .Y(n9892) );
  INVX2TS U13693 ( .A(n9537), .Y(n9538) );
  INVX2TS U13694 ( .A(n11161), .Y(n11162) );
  INVX2TS U13695 ( .A(n11200), .Y(n11201) );
  INVX2TS U13696 ( .A(n10063), .Y(n10064) );
  INVX2TS U13697 ( .A(n10725), .Y(n10726) );
  INVX2TS U13698 ( .A(n10339), .Y(n10341) );
  INVX2TS U13699 ( .A(n9461), .Y(n9462) );
  INVX2TS U13700 ( .A(n11167), .Y(n11169) );
  CLKINVX2TS U13701 ( .A(n12738), .Y(n12717) );
  INVX2TS U13702 ( .A(n9529), .Y(n9530) );
  INVX2TS U13703 ( .A(n10027), .Y(n10028) );
  INVX2TS U13704 ( .A(n9365), .Y(n9366) );
  INVX2TS U13705 ( .A(n10334), .Y(n10336) );
  INVX2TS U13706 ( .A(n10703), .Y(n10705) );
  INVX2TS U13707 ( .A(n9525), .Y(n9526) );
  INVX2TS U13708 ( .A(n10353), .Y(n10355) );
  INVX2TS U13709 ( .A(n10317), .Y(n10318) );
  INVX2TS U13710 ( .A(n10047), .Y(n10048) );
  INVX1TS U13711 ( .A(n9350), .Y(n9351) );
  INVX2TS U13712 ( .A(n10330), .Y(n10331) );
  INVX2TS U13713 ( .A(n9361), .Y(n9362) );
  INVX2TS U13714 ( .A(n10087), .Y(n10088) );
  INVX2TS U13715 ( .A(n10720), .Y(n10722) );
  INVX2TS U13716 ( .A(n10091), .Y(n10092) );
  INVX2TS U13717 ( .A(n10043), .Y(n10044) );
  CLKINVX2TS U13718 ( .A(n9843), .Y(n9844) );
  INVX2TS U13719 ( .A(n10358), .Y(n10359) );
  INVX2TS U13720 ( .A(n10095), .Y(n10096) );
  INVX2TS U13721 ( .A(n11179), .Y(n11180) );
  INVX2TS U13722 ( .A(n9369), .Y(n9370) );
  INVX2TS U13723 ( .A(n9851), .Y(n9852) );
  INVX2TS U13724 ( .A(n10353), .Y(n10354) );
  CLKINVX2TS U13725 ( .A(n12737), .Y(n12718) );
  INVX2TS U13726 ( .A(n9354), .Y(n9355) );
  INVX2TS U13727 ( .A(n9373), .Y(n9374) );
  INVX2TS U13728 ( .A(n10317), .Y(n10319) );
  INVX2TS U13729 ( .A(n11195), .Y(n11196) );
  CLKINVX2TS U13730 ( .A(n12738), .Y(n12715) );
  INVX2TS U13731 ( .A(n9819), .Y(n9820) );
  INVX2TS U13732 ( .A(n10751), .Y(n10753) );
  INVX2TS U13733 ( .A(n9895), .Y(n9896) );
  INVX2TS U13734 ( .A(n11161), .Y(n11163) );
  INVX2TS U13735 ( .A(n11200), .Y(n11202) );
  INVX2TS U13736 ( .A(n9285), .Y(n9286) );
  INVX2TS U13737 ( .A(n9450), .Y(n9451) );
  INVX2TS U13738 ( .A(n9533), .Y(n9534) );
  INVX2TS U13739 ( .A(n10708), .Y(n10709) );
  INVX2TS U13740 ( .A(n10736), .Y(n10738) );
  INVX2TS U13741 ( .A(n10334), .Y(n10335) );
  INVX2TS U13742 ( .A(n10746), .Y(n10748) );
  INVX2TS U13743 ( .A(n10039), .Y(n10040) );
  INVX2TS U13744 ( .A(n9347), .Y(n9348) );
  INVX1TS U13745 ( .A(n9344), .Y(n9345) );
  INVX2TS U13746 ( .A(n11189), .Y(n11190) );
  INVX2TS U13747 ( .A(n10358), .Y(n10360) );
  INVX2TS U13748 ( .A(n9521), .Y(n9522) );
  INVX2TS U13749 ( .A(n9453), .Y(n9454) );
  INVX2TS U13750 ( .A(n9827), .Y(n9828) );
  CLKINVX2TS U13751 ( .A(n10708), .Y(n10710) );
  INVX2TS U13752 ( .A(n10339), .Y(n10340) );
  CLKINVX2TS U13753 ( .A(n11195), .Y(n11197) );
  INVX2TS U13754 ( .A(n9795), .Y(n9796) );
  INVX2TS U13755 ( .A(n10344), .Y(n10345) );
  INVX2TS U13756 ( .A(n9281), .Y(n9282) );
  CLKINVX2TS U13757 ( .A(n12738), .Y(n12716) );
  INVX2TS U13758 ( .A(n9811), .Y(n9812) );
  INVX2TS U13759 ( .A(n9879), .Y(n9880) );
  CLKINVX2TS U13760 ( .A(n12737), .Y(n12720) );
  INVX2TS U13761 ( .A(n10363), .Y(n10364) );
  INVX2TS U13762 ( .A(n11167), .Y(n11168) );
  INVX2TS U13763 ( .A(n9446), .Y(n9447) );
  INVX2TS U13764 ( .A(n9855), .Y(n9856) );
  INVX2TS U13765 ( .A(n10348), .Y(n10349) );
  CLKBUFX2TS U13766 ( .A(n12655), .Y(n12606) );
  CLKBUFX2TS U13767 ( .A(n12655), .Y(n12612) );
  CLKBUFX2TS U13768 ( .A(n12655), .Y(n12611) );
  INVX2TS U13769 ( .A(sa21[4]), .Y(n10725) );
  INVX2TS U13770 ( .A(sa02[1]), .Y(n11173) );
  INVX2TS U13771 ( .A(sa02[6]), .Y(n10730) );
  INVX2TS U13772 ( .A(sa33[7]), .Y(n10751) );
  INVX2TS U13773 ( .A(sa33[3]), .Y(n10741) );
  INVX2TS U13774 ( .A(sa23[2]), .Y(n11200) );
  INVX2TS U13775 ( .A(sa33[6]), .Y(n10746) );
  INVX2TS U13776 ( .A(sa10[4]), .Y(n10698) );
  INVX2TS U13777 ( .A(sa13[6]), .Y(n11195) );
  INVX2TS U13778 ( .A(sa30[7]), .Y(n10714) );
  INVX2TS U13779 ( .A(sa22[2]), .Y(n11189) );
  INVX2TS U13780 ( .A(sa13[3]), .Y(n10736) );
  INVX2TS U13781 ( .A(sa30[3]), .Y(n10708) );
  INVX2TS U13782 ( .A(sa12[2]), .Y(n11184) );
  INVX2TS U13783 ( .A(sa02[3]), .Y(n11179) );
  INVX2TS U13784 ( .A(sa00[0]), .Y(n11161) );
  INVX2TS U13785 ( .A(sa01[7]), .Y(n10720) );
  INVX2TS U13786 ( .A(sa11[2]), .Y(n11167) );
  INVX2TS U13787 ( .A(sa20[3]), .Y(n10703) );
  CLKINVX2TS U13788 ( .A(n9594), .Y(n9596) );
  CLKINVX2TS U13789 ( .A(n9314), .Y(n9316) );
  CLKINVX2TS U13790 ( .A(n9614), .Y(n9616) );
  CLKINVX2TS U13791 ( .A(n9609), .Y(n9611) );
  CLKINVX2TS U13792 ( .A(n9336), .Y(n9338) );
  CLKINVX2TS U13793 ( .A(n9599), .Y(n9601) );
  CLKINVX2TS U13794 ( .A(n9464), .Y(n9466) );
  CLKINVX2TS U13795 ( .A(n9319), .Y(n9321) );
  CLKINVX2TS U13796 ( .A(n9404), .Y(n9406) );
  CLKINVX2TS U13797 ( .A(n9478), .Y(n9480) );
  CLKINVX2TS U13798 ( .A(n9562), .Y(n9564) );
  CLKINVX2TS U13799 ( .A(n9619), .Y(n9621) );
  CLKINVX1TS U13800 ( .A(w3[27]), .Y(n9599) );
  CLKINVX1TS U13801 ( .A(w3[29]), .Y(n9609) );
  CLKINVX1TS U13802 ( .A(w3[26]), .Y(n9594) );
  CLKINVX1TS U13803 ( .A(w3[9]), .Y(n9562) );
  CLKINVX1TS U13804 ( .A(w1[17]), .Y(n9404) );
  CLKINVX1TS U13805 ( .A(w2[1]), .Y(n9464) );
  CLKINVX1TS U13806 ( .A(w3[31]), .Y(n9619) );
  INVXLTS U13807 ( .A(w2[11]), .Y(n9483) );
  INVXLTS U13808 ( .A(w3[3]), .Y(n9553) );
  INVXLTS U13809 ( .A(n2353), .Y(n10538) );
  INVXLTS U13810 ( .A(n2286), .Y(n10564) );
  INVXLTS U13811 ( .A(n1727), .Y(n11136) );
  INVXLTS U13812 ( .A(n5309), .Y(n11208) );
  INVXLTS U13813 ( .A(n5394), .Y(n11223) );
  INVXLTS U13814 ( .A(n3557), .Y(n11406) );
  INVXLTS U13815 ( .A(n2329), .Y(n11490) );
  INVXLTS U13816 ( .A(n3625), .Y(n12045) );
  INVXLTS U13817 ( .A(n3554), .Y(n12253) );
  AOI32XLTS U13818 ( .A0(n10314), .A1(n9175), .A2(n4334), .B0(n12200), .B1(
        n11769), .Y(n4332) );
  AOI22XLTS U13819 ( .A0(n12145), .A1(n10644), .B0(n12372), .B1(n11490), .Y(
        n2888) );
  AOI22XLTS U13820 ( .A0(n11489), .A1(n12139), .B0(n12373), .B1(n11110), .Y(
        n2328) );
  AOI22XLTS U13821 ( .A0(n12132), .A1(n10637), .B0(n12368), .B1(n11494), .Y(
        n2812) );
  AOI22XLTS U13822 ( .A0(n11495), .A1(n12124), .B0(n12366), .B1(n11094), .Y(
        n2261) );
  AOI31XLTS U13823 ( .A0(n9286), .A1(n11461), .A2(n10001), .B0(n7928), .Y(
        n7922) );
  AOI22XLTS U13824 ( .A0(n11422), .A1(n11512), .B0(n10679), .B1(n11519), .Y(
        n3107) );
  AOI21XLTS U13825 ( .A0(n4475), .A1(n10318), .B0(n11779), .Y(n4297) );
  OAI21XLTS U13826 ( .A0(n10520), .A1(n12451), .B0(n10967), .Y(n2482) );
  AOI22XLTS U13827 ( .A0(n12373), .A1(n11489), .B0(n11845), .B1(n10644), .Y(
        n2675) );
  AOI31XLTS U13828 ( .A0(sa21[4]), .A1(n2940), .A2(n11846), .B0(n2941), .Y(
        n2934) );
  AOI22XLTS U13829 ( .A0(n12138), .A1(n11845), .B0(n11937), .B1(n2409), .Y(
        n2406) );
  AOI31XLTS U13830 ( .A0(n10699), .A1(n2864), .A2(n11839), .B0(n2865), .Y(
        n2858) );
  AOI221XLTS U13831 ( .A0(n11247), .A1(n12505), .B0(n11270), .B1(n11209), .C0(
        n6421), .Y(n6399) );
  AOI22XLTS U13832 ( .A0(n10864), .A1(n12503), .B0(n10995), .B1(n12264), .Y(
        n6199) );
  AOI211XLTS U13833 ( .A0(n12503), .A1(n10994), .B0(n5454), .C0(n6418), .Y(
        n6773) );
  AOI221XLTS U13834 ( .A0(n11310), .A1(n12509), .B0(n11284), .B1(n11392), .C0(
        n4693), .Y(n4671) );
  AOI22XLTS U13835 ( .A0(n10888), .A1(n12507), .B0(n10773), .B1(n12216), .Y(
        n4436) );
  AOI211XLTS U13836 ( .A0(n12509), .A1(n10772), .B0(n3765), .C0(n4690), .Y(
        n5032) );
  AOI221XLTS U13837 ( .A0(n11295), .A1(n12521), .B0(n11318), .B1(n11221), .C0(
        n6493), .Y(n6471) );
  AOI22XLTS U13838 ( .A0(n10880), .A1(n12519), .B0(n11007), .B1(n12273), .Y(
        n6239) );
  AOI211XLTS U13839 ( .A0(n12518), .A1(n11006), .B0(n5520), .C0(n6490), .Y(
        n6831) );
  AOI221XLTS U13840 ( .A0(n11358), .A1(n12525), .B0(n11333), .B1(n11404), .C0(
        n4621), .Y(n4599) );
  AOI22XLTS U13841 ( .A0(n10905), .A1(n12524), .B0(n10761), .B1(n12223), .Y(
        n4396) );
  AOI211XLTS U13842 ( .A0(n12523), .A1(n10760), .B0(n3699), .C0(n4618), .Y(
        n4974) );
  AOI22XLTS U13843 ( .A0(n12499), .A1(n12213), .B0(n11286), .B1(n3594), .Y(
        n3883) );
  AOI22XLTS U13844 ( .A0(n10116), .A1(n3671), .B0(n10415), .B1(n12016), .Y(
        n4314) );
  AOI31XLTS U13845 ( .A0(sa00[2]), .A1(n3947), .A2(n12017), .B0(n3948), .Y(
        n3946) );
  AOI211XLTS U13846 ( .A0(n3925), .A1(n12018), .B0(n4566), .C0(n4567), .Y(
        n4565) );
  AOI22XLTS U13847 ( .A0(n11218), .A1(n10429), .B0(n9934), .B1(n12045), .Y(
        n4241) );
  AOI22XLTS U13848 ( .A0(n10853), .A1(n6089), .B0(n10863), .B1(n12234), .Y(
        n6082) );
  AOI22XLTS U13849 ( .A0(n10899), .A1(n4223), .B0(n10887), .B1(n12231), .Y(
        n4216) );
  AOI31XLTS U13850 ( .A0(n4086), .A1(n9144), .A2(n12420), .B0(n4683), .Y(n4676) );
  AOI22XLTS U13851 ( .A0(n12498), .A1(n9638), .B0(n12419), .B1(n11393), .Y(
        n4437) );
  AOI22XLTS U13852 ( .A0(n12501), .A1(n12421), .B0(n9643), .B1(n9114), .Y(
        n4115) );
  AOI31XLTS U13853 ( .A0(n5830), .A1(n9430), .A2(n12392), .B0(n6411), .Y(n6404) );
  AOI22XLTS U13854 ( .A0(n12513), .A1(n5875), .B0(n12391), .B1(n11210), .Y(
        n6200) );
  AOI22XLTS U13855 ( .A0(n12510), .A1(n12393), .B0(n9731), .B1(n9297), .Y(
        n5859) );
  AOI31XLTS U13856 ( .A0(n4030), .A1(n9347), .A2(n12436), .B0(n4611), .Y(n4604) );
  AOI22XLTS U13857 ( .A0(n12514), .A1(n4075), .B0(n12435), .B1(n11406), .Y(
        n4397) );
  AOI22XLTS U13858 ( .A0(n12516), .A1(n12437), .B0(n9647), .B1(n9107), .Y(
        n4059) );
  AOI31XLTS U13859 ( .A0(n5886), .A1(n9343), .A2(n12408), .B0(n6483), .Y(n6476) );
  AOI22XLTS U13860 ( .A0(n12529), .A1(n12591), .B0(n12407), .B1(n11223), .Y(
        n6240) );
  AOI22XLTS U13861 ( .A0(n12527), .A1(n12409), .B0(n9735), .B1(n9307), .Y(
        n5915) );
  INVXLTS U13862 ( .A(rst), .Y(n12654) );
  NOR4X1TS U13863 ( .A(n7773), .B(n7200), .C(n7907), .D(n7908), .Y(n6984) );
  CLKBUFX2TS U13864 ( .A(n1336), .Y(n12660) );
  CLKBUFX2TS U13865 ( .A(n1276), .Y(n12661) );
  CLKBUFX2TS U13866 ( .A(n1271), .Y(n12662) );
  CLKBUFX2TS U13867 ( .A(n1292), .Y(n12663) );
  CLKBUFX2TS U13868 ( .A(n5204), .Y(n12664) );
  CLKBUFX2TS U13869 ( .A(n3407), .Y(n12665) );
  CLKBUFX2TS U13870 ( .A(n1438), .Y(n12666) );
  CLKBUFX2TS U13871 ( .A(dcnt[0]), .Y(n12667) );
  INVX2TS U13872 ( .A(n3364), .Y(n12668) );
  AOI22XLTS U13873 ( .A0(n3363), .A1(n3364), .B0(n1629), .B1(n1784), .Y(n3362)
         );
  INVXLTS U13874 ( .A(n5247), .Y(n12669) );
  CLKBUFX2TS U13875 ( .A(n3339), .Y(n12670) );
  CLKBUFX2TS U13876 ( .A(sa00[1]), .Y(n12671) );
  CLKBUFX2TS U13877 ( .A(n1317), .Y(n12672) );
  CLKBUFX2TS U13878 ( .A(n5126), .Y(n12673) );
  CLKBUFX2TS U13879 ( .A(n3332), .Y(n12674) );
  AOI22XLTS U13880 ( .A0(n3330), .A1(n9073), .B0(n3332), .B1(n9130), .Y(n3328)
         );
  CLKBUFX2TS U13881 ( .A(n5150), .Y(n12675) );
  CLKBUFX2TS U13882 ( .A(n3353), .Y(n12676) );
  CLKBUFX2TS U13883 ( .A(n1358), .Y(n12677) );
  CLKBUFX2TS U13884 ( .A(n6953), .Y(n12678) );
  INVX2TS U13885 ( .A(n2558), .Y(n12679) );
  CLKBUFX2TS U13886 ( .A(sa01[6]), .Y(n12680) );
  INVX2TS U13887 ( .A(n6352), .Y(n12681) );
  AOI22XLTS U13888 ( .A0(n6990), .A1(n6924), .B0(n9156), .B1(n1566), .Y(n7032)
         );
  AOI22XLTS U13889 ( .A0(n6932), .A1(n6933), .B0(n1608), .B1(n1644), .Y(n6931)
         );
  AOI22XLTS U13890 ( .A0(n3337), .A1(n3338), .B0(n9134), .B1(n1996), .Y(n3336)
         );
  NOR3BX1TS U13891 ( .AN(sa00[0]), .B(n9236), .C(n9208), .Y(n3924) );
  CLKBUFX2TS U13892 ( .A(n12764), .Y(n12762) );
  CLKBUFX2TS U13893 ( .A(n12764), .Y(n12761) );
  CLKBUFX2TS U13894 ( .A(n12759), .Y(n12747) );
  CLKBUFX2TS U13895 ( .A(n12759), .Y(n12748) );
  CLKBUFX2TS U13896 ( .A(n12762), .Y(n12741) );
  CLKBUFX2TS U13897 ( .A(n12760), .Y(n12746) );
  CLKBUFX2TS U13898 ( .A(n12762), .Y(n12744) );
  CLKBUFX2TS U13899 ( .A(n12761), .Y(n12742) );
  CLKBUFX2TS U13900 ( .A(n12760), .Y(n12745) );
  CLKBUFX2TS U13901 ( .A(n12763), .Y(n12760) );
  CLKBUFX2TS U13902 ( .A(n12757), .Y(n12735) );
  CLKBUFX2TS U13903 ( .A(n12762), .Y(n12733) );
  CLKBUFX2TS U13904 ( .A(n12762), .Y(n12734) );
  CLKBUFX2TS U13905 ( .A(n12761), .Y(n12740) );
  CLKBUFX2TS U13906 ( .A(n12758), .Y(n12749) );
  CLKBUFX2TS U13907 ( .A(n12763), .Y(n12758) );
  CLKBUFX2TS U13908 ( .A(n12759), .Y(n12736) );
  CLKBUFX2TS U13909 ( .A(n12763), .Y(n12759) );
  CLKBUFX2TS U13910 ( .A(n12765), .Y(n12763) );
  CLKBUFX2TS U13911 ( .A(n12761), .Y(n12743) );
  CLKBUFX2TS U13912 ( .A(n12761), .Y(n12739) );
  CLKBUFX2TS U13913 ( .A(n12765), .Y(n12764) );
  CLKBUFX2TS U13914 ( .A(n12760), .Y(n12756) );
  INVX2TS U13915 ( .A(n12746), .Y(n12693) );
  INVX2TS U13916 ( .A(n12745), .Y(n12694) );
  INVX2TS U13917 ( .A(n12746), .Y(n12691) );
  INVX2TS U13918 ( .A(n12749), .Y(n12684) );
  INVX2TS U13919 ( .A(n12748), .Y(n12686) );
  INVX2TS U13920 ( .A(n12747), .Y(n12690) );
  INVX2TS U13921 ( .A(n12747), .Y(n12689) );
  INVX2TS U13922 ( .A(n12748), .Y(n12687) );
  INVX2TS U13923 ( .A(n12747), .Y(n12688) );
  INVX2TS U13924 ( .A(n12748), .Y(n12685) );
  INVX2TS U13925 ( .A(n12746), .Y(n12692) );
  CLKBUFX2TS U13926 ( .A(n12765), .Y(n12757) );
  INVX2TS U13927 ( .A(n12749), .Y(n12683) );
  INVX2TS U13928 ( .A(n12749), .Y(n12682) );
  CLKBUFX2TS U13929 ( .A(n9039), .Y(n12738) );
  CLKBUFX2TS U13930 ( .A(n12765), .Y(n12737) );
  CLKBUFX2TS U13931 ( .A(n12759), .Y(n12755) );
  CLKBUFX2TS U13932 ( .A(n9039), .Y(n12753) );
  CLKBUFX2TS U13933 ( .A(n9039), .Y(n12752) );
  CLKBUFX2TS U13934 ( .A(n12757), .Y(n12750) );
  CLKBUFX2TS U13935 ( .A(n12757), .Y(n12751) );
  CLKBUFX2TS U13936 ( .A(n12756), .Y(n12754) );
  NOR2BX1TS U13937 ( .AN(n9059), .B(n9071), .Y(n2469) );
  NAND3BX1TS U13938 ( .AN(n11162), .B(n9204), .C(n9208), .Y(n3954) );
  NOR2BX1TS U13939 ( .AN(n8648), .B(n9617), .Y(n7155) );
endmodule

