library verilog;
use verilog.vl_types.all;
entity wddl_or_tb is
end wddl_or_tb;
