module not (a_i, out );
  input a_i;
  output out;

INVXLTS U0 ( .A(a_i), .Y(out) );

endmodule
