*include model and subckts
.lib '/tools2/courses/ee6321/share/IBM_PDK/cmrf8sf/relDM/HSPICE/models/allModels.inc' tt
.include '/tools2/courses/ee6321/share/IBM_PDK/cmrf8sf/relDM/HSPICE/models/design.inc'
.include '/user4/spring13/jy2525/lib/subckts.sp'


.TEMP 25
*define options
 .option post=1
 .option accurate=1
 .option gmin=1e-15
 .option gmindc=1.0e-15
 .option method=gear

*circuit instantiation
x1DFFTRX2TS clk d q nett_0 reset gnd vdd DFFTRX2TS
x2DFFTRX2TS clk nd qb nett_1 reset gnd vdd DFFTRX2TS
x3DFFTRX2TS clk q q1 nett_2 reset gnd vdd DFFTRX2TS
x4DFFTRX2TS clk qb q2 nett_3 reset gnd vdd DFFTRX2TS

x2INVXLTS nd d gnd vdd INVXLTS

*power and input signals
vclk clk 0 PULSE(0.01 1.2 0 100n 100n 1u 2u)
vd d 0 PULSE(0.01 1.2 0 100n 100n 2u 4u)
vreset reset 0 dc=1.2   
vgnd gnd 0 dc=0
vwddlffvdd vdd 0 dc=1.2

*measurements
.TRAN 300n 10u
.PLOT TRAN P(vwddlffvdd)
.end

