OR2XLTS U0 ( .A(a_i), .B(b_i), .Y(out) );
endmodule