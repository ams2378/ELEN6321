INVXLTS U0 ( .A(a_i), .Y(out) );
endmodule