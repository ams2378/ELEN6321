.TEMP 25
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2

xu4 n6 n7 gnd vdd INVX1TS
.END
