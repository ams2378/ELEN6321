library verilog;
use verilog.vl_types.all;
entity wddland_tb is
end wddland_tb;
