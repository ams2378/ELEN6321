.TEMP 25
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2

xu8 a_i b_i n5 gnd vdd AND2XLTS
.END
